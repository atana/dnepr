XlxV38EB    1e64     672�u=���������qbT���9�S�����%IgrB�=��_�<�j�)���i��C�pgl�e=��HјW8�o`ܳ9A��{w{z$ڌ���Bǌ����%�Th��-����r	vM���Ba�>�D�[e�m����b��J�������H~��ƕy��a&�FW��!oGX?`1��o�&��VB�ݥ9x�N�,.
�˓8������%��Ʒ��)B�[`����@���D W�N\0�]���2�#�WQ6�߈�@����o�TRJ�:��9��D��l����Ԥ��ɘP�? GG�R�;w�貒�&Z;P69�G�.�J��i˷�[ͨ,�-x1O�Qd,�!4�g5��S���X8�sT�X�
�;����W<�����9�շ#;�|���t��a�:�_�!>��P��>qg�i���P5]�*���
�Ȼb�i%�r����:��`?�)w��N0��q���{f��"��u�oMW�Qӎ-l����5]I(��۳��)��&�ǽn�嶐PS��ČW�+����Z���e��t=��h�ҎX%�q �e�Hi0E��[N�`���	RB��-~�t~,Ff8�8�J�Z��*~-�;�]�)��������ܴ�C#���L�yW �����ax<H�[9�i��GAy��0�n��Ҿ�G�m��Zr>�@��\Q��W��u1�	"����H���.��"����լJ�/p-��K���;�6P�����w{}���/�z��s/W$��]���/-�G~�;֚���3{T�����<�Ǖ�(�Fq�,��&AU8Y9��P��Ү��A�wh6��v0��7ݫ&�Ú���k�#p*�p���r�l�!<�+T*��*���M�O����i>�\����Z~����#������ޑ����$�M3�uD�$�����k 1�Κ�l%�O����4f�_�����1s���Y-_('�IG�����0�9P����ĉ��mv�ש�|�t�SR��T~7�t�e�8��0~j����\suuıw�$x&0/�Z��~ѯύY��_Z������K�X��<]�-�;��a�����!�w�Ŗw��)�!�Œ_a� A�Í���Cz�
�������榸ܣ V�,AY���y۽��9���F�Ӵlm��ZwMsHz5r��;CH�S�����6}%�!'Jߩ���23g{=��S}8����ĸ<,��Թ$�fR����!��(k҄�4�̀@�1�-�*�B�E�2U	U�+�~��0�I�L�(���C��`���������h\4��ףCL{uk�l|/���_�k`Ύ�&��B�ʮ5ѷh'�E�'��N�䋘n~�h��a+ɟ��O� lX*�Rv5�%j��7Ä�iz�2pҋ҇��vci��o��12¾��	7�-��]ӳj!�@D�����4�u�1�h��y�*�6�q�L]5�1���:�p�.,TC�	��ג��L9\ǋDʭ_к$�.\�t��cQ��Pl�0��*=�j��_� �0l�Av�����[`� �ݡ�3j^��u����B6��s'�8��A�,Zn�Wz`x�(ބ��'w�������H�