XlxV38EB    143d     501zH�H;��g� ſo>V�R���F�hK�yf ]�pP�x3�������|�0�-Z��Z�+�wڌ��t�6�A+�_;��3m��mM;�?ྴ&DU�5)�L,&	�_!�J�� ��Ǒ��es��0����D�C�.-X�l�i�,�8�aLe�:�1��n�#�]�.�2¡D�'H�4f��lgtpB�g[�Ñ���j0�F������cN����/��w=?<;!5���x`&���E\��ԞQ�Y#���)����ˬ�ťa�K.��ɾ|�,A��?��5ҳ��m)A`���X:��X{)�.�G$c���� #��e�ƺR��$kbR������z�S�3w�9�N�����I����ƿ'��3q"�����6��~�2l��PV�;�O51��=�#hK`y�}YǴ��J^����L"�м��pP:�����&����EU5)�H%��mw�F��g	�;X�x��
�=r��8k��H�Z'�P��)�!4(^[!�5_���'�9h�w�`:O�����@3�����������Pܯ���;�9 �kۑj��*�3,k���B*a�/�kq4{�[mHl&�܃��yL��5j$˸?�Z�zp�E+�󴷩aM-�|�c�b&�Z	�p���c
�?]��2K_Lf��l�<�&�����c_�c�s\��]��٫|�����|��r�\^�����쳁�?��'j+��x2����K��J����Bc�~�^b׶�&K��MKU�0xW��]�~/,��~�Mϟa];u����z�%��a3�9�n��S֗�&����L���\������X-�2��(������ɗ��{�^��H����A�Q��4�����dt�R��̲��\��	Pg�$�ى�73�)�*Ȑ��ȷ!_h\�k��x��fd)��JRdՈ��r�N�qv����3X���τ��e0��7�� ̤��A��vND�xi���P�E��؅����x5�i�*V�zF�<ڔ�h�N�X����*c���1�)�P��K11Ų=��q:��5Ǝ����B�s%:-�ᦣe"|E ��C��L���0#�=z�Z�TW�\>�;�'��?��E�����E�UEs��	Xh��9��X����C�J�=k��PZ6� �!�j��p"���вL�#�	�&\�T]W�/��ffZ�OT5��G��f�1����]��B �(L�=s�f�}a�=ʱ9s��I�`#�g=��kGT��