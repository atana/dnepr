XlxV38EB    f536    2274 >eIj�NVo�'��W��X@��M��H�w�o�偦6Cu��pC'�W~�mI��/C��k�,-�)��ڧ��"`v��sߍ�)�E�>��B�E?�@�����y-x9Ν��ú�i\�:@;��DО��l�dXB��&��G�dͣI���ѻr��S;K����~�F?χv��ЈKvTf���0���c���.ܷ�y���c$�o6	PQ�*�eM�Yve~�H,� ��r8#���P�@VN��A�`�el��O�W7��(���b1(p�����R`�c�r{���H��V%�k�d��XD�$5�=�-��lL���EU�1�q#c�L^L�z[.hȶh�j䩑���U�?B�=�:�'ROq�jǖ�Er��cƈCy�PK�tp2���C�V�<
Ɩ�&���0-�(�X/N!r��"��;\��B+��4n��)�\y5����R0`X���H>/��H�SsI��1Kr� d�Y��쾸}���1L��6�������j�C�h3��!���	$��T\�>��]ʓ�NF��+�z]KSh��ʟl��I�kKvK�⨯�4�2��*D�[Nۮ@Z�M;�l�t���HE��.�=���x����̼2T�H�S��tpɜ'1�G�W	pl�o��-�G�u�gc_��8����)���AzI�ֆ�{��.�'^&sˉ�68�i�N�2�LbE��G�����r��#V�Z٥�w�|� Cs� Ҏ��R�|���u����4v���q��ߖ��e������t���}׉QO��.RX�E<wG��n�	G1�	��RN3��Fdz���|��X��	9J���ΧĨby��}�,�� �w�r�����)T��!@[��y��~�f�W��S��|�����M��kQ�!���C@(i�4�0�BeAT���c�k8�-eX�:@�F����&eZ�8V��[-��p�R�a\�RR��75'�9�ao.����%$�3Y�{��f�{�^�=nMʰ�~}[�٣#�/�{M�w���Owv��HEI�ks¸ZwRd��%˂(��J�@�`���XE�CXs��j�^\�5Y��i[|�x$V%�������Yi�CV�+UE�.��k/b��	�BR��l�X*E�G��!xo3�g����-w
֐r4/����f^���1.�T�L�OQ�,eT�Æ�k#u3O��ˊ�ء\�v�2���M;�L]�顽Q&�Cv?!� ���RI�c���bo�Qu���X�>���EX!i����U��jL�c �����ʇy���7+��4@46�]�����f��ў���!�S���-�Ob�T���{	�^�0���o��Q�cd��E���-d�(eX���ʒ;}�¦�=;��N'��OV�������l1�\ n��^�p�ι�<w��V�M�P������[#�˸ۯ0����ܸX�x_C"�4�2�=�m����,�ψ~ʌ�L!����'�� ����a���T�q���&1�!b�29k���ltѼD!x�7�G蒫Ft�p�����M�,ǎ�A	�H�%H8o��QSEݏc��B�q%�b�9���/>+-l�,�M��c����Z˔O��o�|�0�)�������·���V0��~��:����0��G��ڱ"�*jlI���Pkx��$n�f�N���Q��?��3�6'A��:��,����10�qMG��|=�:������n���{�i|l�qҤ�g��s4��n��~	�'�E�֪��L��7H���&Dt�J׊%
���O[�9*e۩[���(J��FW�j
sΦ""T;����R=���O	�EM@��𤳟�sS�B����� 	�ԯ��"M��u*��L͎Q&�����M���t&`�f��\�6~�3����u҃�Z�gh��o�4�i�	�sAS�[���XR�Z_n��Y@�bv��G�&����t�i4>B��(N�}6<>n�m�������E��	R$&)��Q��]�34����yn~j��r����r�#m��h�"P֝vٌ�Mr�C\��Yzv��kG*��6��bW#g��EdA�=���*����N2���_�@�$�#Cp�`p���N)���{$!�喃Ԟ������
�޸�wt�ZX%����1xq������C*�|��9��S��m��v8��9΄#+8�j�w�+�ZG.h��K�6D��ëU��"�`�V�RX���	�R�$䨓Ȓy��r(����J��oE�Z���,�=2��NA�-e���ЋY��.�5��À��O�ߘ�j�����"�;^���C��D���Z����B������w'�7,=bAt��2A���IΣ���y�p_ 4������m7��5��z�d__��&,������I���D�*�et���;�n��<�T����E�/A��K5��{	���-y\}��G��K��Jc�Me���W���0	�2|3
�zl�l\�ǁ�ݗ$�OXY��6�
��kh�=�w�����a�ט��sP�;�U���y�|�`?W*\v{H��]Ϸ�]t�=��踭����Ip�B�а�x��������֎I9$���L!e8���؝�N�Q���9��l�=Dǳ�rڭ:���X6�[��!�׸��a�����~�H:[O�vv��Qڎ}E�e>絺��H�Wj�r����BB�Jp�d\���;~2
ϒ0{r>��0�qR�bt�g��1��_A}h�߬I�۱�/u���	��H����x��Z��7�ko_o�QH���6#�<�40KE�����������҅�e%~}^�&�<ׯ��$�
����]��)��c���h��@��ME"us�pȈ�^�3ڢ���4����;Ǩ�)�L~)�][��2(�w����,��K�	�������~g��E�1�1��Z�U'��@kK��.�V���\R�$�Aଫ$�2����!x`���w,�_��]�U�=�R�s���ll���5ͮr�{	sE "�����Vƽ��b*�"
��[oJ�E�A��X�������WΎQa�L\Ђ�%�c%�/�Z���a^�/�����$��}��:��px&f��ahX�l���u�[(s�uѣD_��9�.�/���\1�����ظ�?+�O�'6*���^�o[�rl108�!�y��7�l3S]pծ�-����{����(s7�A5D��m6�̴�L����M�ں d{��>��ѹ�s��Tab�B�s��p�K�*E�kء��87�r�r��k�8��r��4pJ�#R-:4CkD;Ź?P˛Pf���nLqAu��(L�6�����y]���m%P$�%����Y�Fti�!�K����QH�m_��EC��k9�U�dly� ^�T�wmS�Y΀�IF( {�b�e�_�[���iG�>�RW�A_��x��#O��D�+�d��Wx?QX���t�U�B�4��𫲛#����f�ǎ��^�xw���V�I@e������/�8���$�OE��|�Z|Vߗ�D�xx�{6aa1a^�S���%���Qs��7?Y2j�ԃ[��h������<�6��q#~��c��i
����A�%-<�yӄh�Dȼز+}�o*�Gm�0k�Ǥ�����꼓�5�+�f����V5���y�r��j"�d)O��?D/�y]1���q�r��q�R��u�_��J;@�����P����x����2�~��ȃON����������~�ǰX���&�����-�O�7��W��'�2�%5D���vn�b���Z�
pWUZ�M��{֢�Cxb�u1��A�	נ�Xt�䎚W�?]�+a�:4�����Fc��wi.Z�`��)�{��86q���N�7�F����+&��Wz���m5���hae���$��0���:gn׷�N��^<�C��ZʾwԊz��Nej�o�SB2���J�,Qyz��R}z2s�R^�
�Ƥ^uyKO�*Q��}}l_�^c\���+>�H�'m�-d��V������κ�(����YI{�|b'�KY�z�3߀�'(1�"����*�I�xq6�>*�L/-���#̄g�/�� �86�ߕf�f��|���Ӊ�4������q~�8�GLPE�< �ԡ�8�IM�]�L9�}��7zE?5����5���p�j�W
�`c�3���ɮ��&&􏚃&�c��G�i$����Xͤ��e�H��A��īܒz�l?���CBE�\Q�$�����{�[�6�?��e�O�h���1����b-��t�Ϛ^��"���yBY�m�������Z	�a�,�(���_�q*x���U
��q��ڬ�L�c����LkE�.��:��}%'���9�I�Emfu���,����z�k-�Bm��VA��A.K�>����F_�����_�8u�QǖDޱP���W��+d�5�)Et�V�j�	��H��	o�B��c9���T�c?���m�X:J��R��qFM��1T����kDr*�-[Xr�?�v�>\p�,p7ޱ�������DH�+Ỗ_A��kt��b51��̾��4�d�����e�@8���륒%��n�*_'<�m̊:Â�X<�Ч.;U>�ix�cGO���z�v�Ih}i%i���e[��Y2��]��m*B`���4A��@������l��ʯ�Ɉ(�]Y������g]	���EN����9Z�����9�mD���偒�/� *��1�@����i����u豤M���r��N/_���5'�+h���ذς�c�M�>,�������7����8�o�_3W�m28��(�7D���nΩ|;A4xv3d�t���J���fa��ت.�~/��́��H§�'��|��'f�S8�HE���J׳#<L8�C�X��rH�1&���p]䳅gYq�W�g���F��}�c�u:��=p��0c�D��I#���(_��ܭ~�6��ʞ��՛�`@I���i�U����o74��G7 ��t՞�1s���>��<��������yp����
n��Y�������l;tO�B+U3�zw�.���#�P���q�����;=�4Y|��"�7v���u��.X���$I�}aC-(����G7F���Ŝ���ܮ�)��KD�ʾ����C	<ƮҼ\7Z�t���]*̫�|FS��@ 8H��	(�|�D��	j��׽��7���Z53`�M'xI�u��n�\Z�'���{�#���K=cN�^�+}wg���
�i�1&U�i�U�t���"���Tqn
��������c|��[��k�Ц�ɖ���&R�_��c��/jL �_7�>�\2�X�۶`�����)S��$Z
�c�v��Cw�6�E���?2?Ԕ����ʵ��˽T8wڍ�1MjQ����"Y�"k	%��4w���y���U�����* �Lt��I�t��c�i�cZ~u�]Ӧ±Y_�(z��=2m����X�Z���ӾJ$J�{��JJ-ȋ���c�"���\����ĺV�Izΐ����{d^>�st(rJ��L)ɻT����mp����F��14Vea��2��(ԋ���r�S�V��e���#���Hr��O ��c!,3UD�o���v��9�Vī�����*���b�n�g�'�{-N�q#K;3�6���=ar��k �;�I`6�� s)S]^h���V�;��9��ˢ�ܗ�� m)�భ:8&������73���u{l�r�y�"�5in�<���@��� �c9tY;�ƥ�L�A����DdPԀ��1n@�{(5���Y�ƅXF�1ET�R����T�l��a���o���=�?ڊ��w�D ��ՊS�����4@u^c/�b�,*33���y8".��L��3�E�I������#���f�|>���\v�JJ��|�l�g�Q_�~�돳�	�7�u�@�B"G���+�b�2St��Y�m�_Z��ۈ���4[����/��u�ta�C1��wG�f�K�!�%fp�&6k�]D��/����2�S��p��i�Y�����)��VXjV�Oo���z�k܎����LR�(�k����`�T|�pز?���t�p7yԭo=�x��ܿh�5����`�v��C��[���������(ó����_�c�����ӵx+SL5���ne5]�!��_J�B6�]��_��|��,�k��a���B�1���#��/�vbZ?T�ʲ��d����y���n��V|}z"��s�u��L�s�qDҐEl�y@*��'1��K�[?�au�W?�$�4u������3�(D�V�:F�[�Q*�L�(��CR�4�s2o�9�׸��㹒y�d���ʈ��غq�{��,�<����x��;���P=�$2�#:z'orr`ȎC]f�Z���pr��<��,�W���n��$9@x
��2�����u�S|��Q/��l�ut�:���?��3����Ԇ��,��uC]��:-j��af�����r��W �#X���������A�}���)`P=���`θh�7`I�AO@���.��Q��0Q˦��a�N5�������Sm�w�vy��0���C�{�X�c�e�G��${��b[�#>Y���1`ػ����2n�$����ks�a?�Z7F��nW�0Tw��0o���_���4���8<�����Q�"��F�J5so�
�@�2���Z����x޶��D�l�!m����!ks^*�d��:KN��$���;�5��e+��6%�(#����6m�����)��+z���"�jfLzg���N����H9V���Xl1�&�mj�%���j;������ރS�=�����=�+�M�2 �~�>eZy�BCa�'�쎠/��.AT�T
)# ��
L,s21A�NEU,��-��nr�I��HQ5[��X���#�x�Ό�|�݉�*n��Q�<z�ri��)�M�d&�lhy,��u9�ׄx�ƨ���p��y>6E�T����~~$�ܲ�ӛ�Qb�G<�3�Ž�]�`0�d��Hj^F�wg���������O��I��;�b�Jw�q�3|WrQ�8�^D�,1q������+*z�H��F�aҍ�c*���e؏</��w��Z"����R+|��'���|�3>�K�MgNY�{_�����V��ì6�Ok�HQ�MȂ
�R��ntw��ƍe��1PA�Kv���)?��C���t������YvM`s�D�qn�'I��@�o�ޙ���aI˻`���?����g�����^�R2�3��&w8��Ibe�~'��&�4������_��a�ؾ�#��?x?�4��ا�)�פh2�̍����n�(?�]H�'8��f�' �ƒ���tB��iL�6�v�f�0�n��$,���V/��R~ͱ���V�O�,[���c�0S;��M,S���I�3�����2%��{�w�YS(}�]��/��Hf�MX�.�������_4�ϕ�N���^� ��r+:�I�9~-gA�Q��ͱ��,ifgX�(o��Y����QY֯�}�B8L/� ��-����x՞����p$�Լ�}�d),�/�M׀����|f�i�lpi�f�R�|�%}������;���ʕ�ӶR�S�gU\��.� 0���B.�4ᱍ�۹�i��t�fnӻ�<��9SM����ױ��.8AkJI`���
�]��p��b<�B�����"��/ͣ?8@�gD$�Y����o��#5�%���θ�����]�����|!�{x_n͑�t뒀�#9<�KIbW`���	|�3뼳B��j��9^��s�7و`�{��yvǅ��E44y��n%�8e�ꛆ���:ϖe��@)���Q��X�5��
��>�i{���$aQ3F�o8��0�'��N���w�F}s�/��>����\<'*�+�&��ILs,���*�>���B}j]z��%4ӹWA㭴8�g	���� .�NN���2j�k��������ku�A���R��* ��k�Yy:��0����R��2*�pIl�&�@�l�|0~M�(㔤� �������˔w���.��Ì��BP<0<d����V�w���=/���/��&�+yH7]s�����VHz٫�]g�����;�}���_n���b�����G�g%�f4S;1S~���S�dp�c�H�޳�U�E���z^e@�T8�+�*�o+�\?��\�n���+`o�@�w[]�N]N���;�d	x
}��4��^ĒɈz����]�H~����om����U��ʨ��<��W��.����
�#N�)
��g��>o�xMD��}��U5�����驼^�p��H�?'���Bi�c9Z�Ey>}7ٝ�����|�p���aP���rAJt������ۚ�'����w�~���\*�:��^m� Ń ��(���CJ)�m+aXv՘s��:^��e|�^��T>�X��W���(MU),�+@-�qʴ����8�O��I"~�U���Q�W������E��!m�����e�@�YF�g�1;.�2:ZѶ]�7]�v�ޖ��c�<��n�*��?��V���<��H�T�]� �P�_�g�!nY%cϮ��s�Ĉ󲣻�Eį ���-�R�f�