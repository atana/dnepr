XlxV38EB    12c7     4d6�E ��6GX�"/�|a��ת���$2d8+���[.,*�m[C�Ʀ8���g&ܜQY8`�
n-z8QCFI"��F8	��ꘊ��S �V�]=�t��X�Nq���Č|�f :v$0XG/1��+�c�-	����,��O����KN�d�Ba�T�����$���0B�kC
F����_@b�2!Z��lY�@J3�n���s�2p�9~�>�5�Cm��-��)܇v������z=Ou `U����C����1W/9Y��x�2�뵭������\�<I� �����>�g2sN��*�o^ =-k���~��oؼ�1o4�F��{�,����Wk�i�m@��8�2 X6�p{p���=8��^�o52uv�j�|�.�/�gܞ�01�4�@*`Z�v��Q^]�]�RUj'�򢟈iiJ'�O�#����}"-M%?�ZS���2�|����e��o}$��p@�"2�}��&}�Qvs���!1�|��F�:�3�����@�N5��PZz��m~
��]?�����B���_ս,�j�$��Y�DJA3M���Z ���q����Tl�����xp9i�Jׁ��Z���rDjuxhI��Qu��$�%���ܛ�	>?+n�4�Y՝z}�����B@��<���>�Ǧ^^�zc�2d�y�y�i�����b��E�^������d����Vm|i��m�����&n�W���A�۬,�1��h��@�R���slQ���F#�g����-��)C>ɠ~�2ԫ*�Yc`��n/_'���{��/%�A�{ȶ�U!ipo���ן?���)/EQ��y��ȴi���7�8ǩW�g��bM㓊���V�߄��Od$=����:ʽ�S7"�?$����6��jW���I�k|WZY{�7�������w]�������h˜�;CL�5c�`�������$)q0A%�:��^��o�Rؒ	r��q!;l=�z���������������_����\ ���"	΂��0�M��������B�a'fy�]�X2�XSO�]�����g$��0k�p��4.�)��a@�`%b����T%�N���2���Uܛ�9J}Jh/�g �9~������2��_L�kA�E��ƺ��; ��i�-aIr���k���Ʈ�@6I���j�ԇCʏ�UcVi��S-I~�V�D������d����h� �	A^�=e�如"�?*B