XlxV38EB    87e9    1c59E��u9S�*�����+^J�̑`���|Ս#r6a����~�zj{����#�d�v8��� ���BE�	OP;!Τ���t���M��2�P%z��(^^�K�okՀ0l��S�'Q/<[D)Y40�S�����Na�Ȥ ��F�F��g�E��e�ٛ�_����@�o=*'���R_)����;Q(?�+Ռ��Y��K[��'?�����&0�1H��X��8HI7-az��}������
�	.!������%��&��S�ф=���m�u`3p4T$�`���Sb>:]��������i"�1�/2����ǈʝ(������$%��ͧ}��Bp~���O�;GY֔��|.��E!E+¸�G�t	:�a���0�&�-��
E�? �iId 	$\j����K�T#��p�'j.�ʳRY_F�K���?��ޗ����Mo�3+sU�\��:��v0�]��՛����{ Zx���L��Xp3Z��)�u㽽��B��zI�W⟿��G�RJu"���Vֻb�'�_;���NW��&9��`��.�f���2��qczgl~����od+�CJ��[َ0�,ܘ�4�]�q̘�B�7)*!��,q ������P�}�8����r*f��td�n�`8}��w=?��K��U�7cV��w%��jX��ۢ���H���z"���f�x��1�Kr�Ĺ��ӝK��[�n!�y���XB��em�?�������ȧ�M�ɕ��Q�� ��Qy"�8]ՙ��cy�:�`}I0@+v�n�_�]�[�ZZ�Z���`Pf�M�J�Չ�Mea�/�?Z@_�}}��ګ��IO� �.iW)�>���k
6�:��<F2��ϡ��h��#���.?R#�AF:���G�Dy�	 ݷ�A��8� �C�x��,������T�ιg��AD�?�|B`�O����q-[qFC#*Sw���J�mRd�&k ���KW��]�6*�fQ�Q�w�d��l�/5�J�Z�F�Ïeӈ����j\���-��+���sـ��+dHIj�#(�:y���-#SL|,��\����K$���N���UJ��B�[�8�冚����p��$�Zp���~�96�S#����ۥD���4(�S��bÚeN΂/WWq�.40�0nB�K���Wr�=|g�$�so�
Cؾ�2�ǟ��>eO���?��z�+��Mؕz��}�pf�\
u}ZS{K0�HLl%R�y$a�Y:�3DF�"�J&���緬_%f��K�����8�Q7���:�x�i|���!�é df��/�ٱ���,�Q��"/��j:���\��S�J�J��AT����$?8j�m�}.ݕ�VV�qP3zv2��A�!ˇG8 �Rj�W"Wũ���i�}Ţ^qq�Uε�����0p�/wTT�M�B��'�o�L��LP�0^���GKD� H`���� �/A[�L'PI,?��tЁ��_g�ʠ��ẵ�� �R���֍�}�e�b2� |��-@H���k�������hy��'�����xoy�����,���<���@B{���բ�xj5��-��O�� �H���@K�v ��E�3��0?+*,���� zD�.�L���QE-O]�%�c�M`_�P�
��zF�H�	Qa#O���8
�b�R�և�(l
c��h�Q$U�6ot~�	ԃ��I��<��zM}9�g6U���
���%r�N�Y���U9�vS��AJl�W|��ǐ@�;|R��Z�?|��
�]���� 5Ls�~P��4K��a��>�#������*#u91E��{$�\~8���~����e+�c!�Ӫn,�C��Q�\ ��`�a�uԖ [P	ʌ7�|	{��U^g�����|_2�d�h\*����A�P$ؾ4]-]a&5�7�!�����|�Gˮ �`Σ>��&�ov����xY�"��8UT0��ρҫDi��J��ӿbGf��`�N�L��'����8�~�t���ݯ��ۢ���~@Ϗ��H��,�7O��ū�=j�&��>.�춀���&��3X�qH)�%N�M�x?�\r�� ��B�ݩbP�Q�j�����ldU����1���J#��δW�Ƽ�k��$D�_	�<c�A �i��"jJ9:�>��3-w>�tf�;�� ����f�DI�"ѓ���u�����>��m�:ؼ��q�Q(���~^���i��3�� �ZH^K�r&��x��q��^���J��c@������T���a�}	��i4WIM/-\a��y���?n?��ԛ���_�o��F�����v�u��]���0������ia
��K�E�y~��`��K�$�����WI�*�<���ճn��c-@�+��S��XI=�����O�P6�R�>V���4.��l%�'�}�ن�&u�$R��<��ҡ-4>�
3<\��ˏ#��(�V�Y�t��9�$��m��Nѡ<҅K������^0�P/����,ӆO�p�
�1�߁�m��r#�e��v�F)+����h�ua-�v�ÜV��Rd�mґݓ�U�_��v�d@3o*m�t1/�7�y�9t,T�w�����7J� �Q�L��K�6Ţ�$����V�Z�IW���De��2�T8[�Pr�tz8 TC�';ܕ6�� �5�U����rf�
$��Q\�S�kMUCgZ8�x�h��h=ޱ� ���(KZi&4L�m�J�)����� y4���1��}/"p��JJ�bJ���/����^��:�l�֟O�7^	p�$�B]���#��n{wsA��-���L����9<I|�%QA��G��_�6?�!z�}��Z�MԳ������㌑�iH�U���D�#�W|ە/�N����Q.�v�=
S��2x��rZ�]o�P��>Ò�tR�1�i*c" h�1��=��[c���J��f�S�I�����	s���2`���"�`��ujN��a��s�g$�5���t�]6Eo5z�O������z"G�A�v����HL2�|��baO��K��V2��lp�a��aL�o|�}Z�ȹ�P�r?�$ `�M½6ۏx�&8*(���E������ē��a��fJ1�����gb������>I���M���3Nj&��AK��4cc�.�O��g�=�a�k9�N�eT�u����lD��ڜ�c�
�hD����N�x�C���=#^� ��	�j�+{�c2uu?3�_��4d����DOK�pF����{�S����t��H�o~ǆWT��Df��Y�Uq�eE(nG�m��J��5N��*0&�^~�f�lb?�Ha���I�k�:B�p�L�%E�Q�ţ�$+�Ws�
��|@` o����@�b��J�*�PH�Mv~H��P���!�S���2_ᵤ5`6,�7��'���9#6��]���\�;^(�(ĳg�i��}JΟ��������M����e$�o���	�2r'\�݆��:�62�Px������i��ǬG����Y~����#b���P�ih���%���F�Hf���9�ØC'N\�o@>�YrTdt!)<�^����
�GA�6�|ȜX:��I�$}k8�[�빬�h�%�Ls���uH�a���۠���D��D{�����f�����<��j��J{�4k��>o#�g ��b��0?�-�V��qT{�j�,��k�+�k6�!j�dʌá�}���]=�B�O*�>�td:�0ҏ�>���_����Z}��܆�3J~��zH��#��J�U�ѥ���Ldt<��q$O��0a�6��Ir&����U�K�q��V�VQ3Y�n�qb�""��.��ֳ�3J��b>��0�L�$3�[)��~̶r=���%>��?�z�=�^&R%9���r�Wb#���n��/߹肝�Y"�:����(�:�U<����Y>���F#�3pɈ�lq�5J���q���sT$%Q�Ugü秿~�+'�.r��?2�[|i��R�R�D����=���A(�&dV	��>�/� |M���-{���^�օ���wj���,򥗚�D�.:X�l�ǝ��IG�h��4��&����֑�9�}����Vn_�~u��s�_��A,*��4f��� �v�B������K[T�W�];����ڳ!{UI|�^oMŰ������5g�=�`fi�̔���P�]�i����������Y̖�?F��@����xx<4�8�Q$ �@p-Y@�E�Zk6���Bd:�+�|��Bg��v��_��I���Xz��aԋ������uL@Mh�U�^,�8���se]�(�} ���&��,W�.no����h�$ �&�1.���"��U��M��f���aS֝Z���"�Zj"�\�$d�s�t�v�C�&ʄ9����t��s��K+� �ՠ��O�\>�5�|���t�5���h�G�_nr��u��ϻ�қ��d�2�c�#������Ν��2ܝ������]�B@�x�d1��n��u��Ѻ�@����nJ��������P������	Y~E�u�+HkMa����"��!�K�DB�K�f;�@�����u3�� ,�tkx�,����щ$��a�헵`�s�)�x��y�lTVηU�s��@�Yke�,P�خ���Wޏ�B�\ڏ#��Ҟ���uydT^�FO��sD�e�wYߴ	ه��˔��>& $����ݵ3��Ɏ����X�w�[1o�g0���^:|~h�X�����e�i9��c�>f�}�����a�G�}��QTC�)�6��]0j��@I6�r(�d�(%��V�����o��lrD3��u�M!����l��'N��w��冷.�t��W?��?%�I�:��f�4�ҒM�{�L����_9�]`#���av�Ҽm��G��=�D&�9�k�qsUN��xL��'�?0ݖ�����0�W�1GV���]k��o@�UQꭙ���˟B����>�M͖�it�X��w������8����b��0�<9;Oh��t�캍�z��p���X���6q)	���_W|�$��(�3a��(�~��q
�k�7�li'�u���;9�R~�	�s#5�Z��D�^��"����T ���
���,���W��QXS���f�٨�x��2�"ʶw����Zv��L�N��Î�L���?���2j?�>$#�/�m����� �٠��S�N�G4��n��j�-��.H��^Ν�n��o���R^��52�('%��9p�	�y=�l�MM�#ܴ�@��w���B	���F*���Qz^�p���6��`�1�5�9�NW4R�f&�3�/�v^���Ps��LJ^ʺ8��gLoV�M�(+���IAN-C�V�'l8� ��1}:�3m�T�MÙ�:r�0��|��$\����m�����S�m���8 ��EM��V1�3��e�!3f�r�=�u�}��P%Q�1�H��j���t�3;9~!^����H^z�B�0�TE�z=/e��-TLM۞@�.S��f	��UF�k��0���`�G$ *�6�BSU��[;��pk31���a6���s��v^�U�S�X��b�1m���]�<���F�\��S���`H���:m|h�{^�+s-�Q�Y~bZ市L�mGZ S��������N�}�v�u�����.�E$��T�n�w�}���9�Bz�iS����X�쾰����k8���LpM�{�cq��'G����^M��a��p��ք�zY��d��^� �ݖ��A��yٽ��3�h���QH)b����2�S�ٹA�=�f�S���U��q�sP�e#E�W��;'�ӧ�i�9K������s���j߻Z�ٷ�m� �9aY�}���g~���@�b����C�iҩoiR?ˮ�u����ܺ�]'�e7�<��b&��H�=������K6�-� ��XR��J�wς��h0�������<
W-U3V:؝��t�����
�O�=Y���̗�4>'	1��o�p��t�+�T_z��b���p���ٌ�W!K㡖��J�)�3;$SʇE���ۗ�KC�1!�� ��`E4�;y��2Pn�\��\��w;�@1�E�%Պ�L���d���'�v暈Y�k��91�q�`'�ɯ+��K�7sمm�w���շ��U��E��'N���o�b�Xş��L.��F�Ir"�1�5��S�06�Y��g�����neb�g��WS]�v��[t���
��=j�x��X�p�k@s����DR�#`��߆R7�a����_q���e$C}��Z��ZF���i��h�f��c!�����"�PįLZ{�{�(����@LH܄Y+���ҏQs�o:[S':D���ś:�ĞKiC@(�l��f� 1ʦ���֣�nA�3�9$&��9G�/3������k�gsQ�K��o�v� �?�۝����%!���nJFc���jjh��SSK9�����_?�x,+.<�[|F����Y��`ߐ���9{#�Иo;7���_0NY�F�&nS�FK��U�����%q}�{eȌJ(�#�Z*aO(��$Q��F�6��z�G��$2n�6�^���C�"�y7�X ��4��Է&=;���L#�zE���&O�~����Z���b����Y=S2-��=��U����~��"�RE�HIf��S�[ ���g\�\G�U��Cȡ����9�WV8���*H�P��X�{^������f��d��gLmqf+�f�.�Խ��Ҷ6)�9ǽ8����"Z��Q;�(�7�ܫ��;��o��L�O��h���M��y���J��-k��jl%=�!������s<?�	qڅ@8|�ic����}�P]���}���儻Àg8Ū���*xf�����Po���b	Z8���YIT�a��uE��K�S��
%�"�����y\%4��2�=2�_��ǜ�����8~�S���f��/xg刼�k㚉m��J�vq��	�~%���Ė��fn6�/����D2ޏ����P���N��R�on�4{����T �ō��P��t':23��L�企�8�I~�������^��{����^*2