XlxV38EB    2800     c5as�'#�LI{E���;�1k�G;�lG�Zي�}C�ȴP��X�ZF�*�.|]"��h�{Za�����@V� �ͽGU���X'1������@s"��y �s3P�GN�m{ɶF1^iS\��Ӟi��J�O�Dî�Kit)��WE��T�o�Qt���08D�h2՜/O�Z���ʻ���%����bNk�<��S��"3`ȴ+�D+�I�x6��Yqo�1x�k5���%��t�a?88��d�� ��%��Y�)�-��I��L�����&=����:L�`�M)�=�S��vzg/�9�qE3���_|W��!��YE�x��.�Zi��_����K�U���)�
s��/Z�O��u0[�՟������(wJ�>�/}��w#d=���h,�jy�W�hCH��ν�y�$T�}��;��M[�Х��byZ���!�	@OG�p��H[1Ӯ.=-ʭjG�5���R�8��-YK`���yTN�
q!��"����p�e9���S��3�q�j3)q�(�4	��0V��?௨�֪ȳ5��TZ(��'����<_�!�{kx(_x��SQ�z���s�$y�alI���[&jY��l���0	�T�y���z�#?��ȃ?�E�@}�)�� Lv���6U��Z�̒8E��OY��l�i����Ȳ�h\�g�d�M�Jm��c_�v�^���JUc�MR��h��Xx��n!N��E�D�r?��Tu���(j���Z��p�l�"%8��I�`@����Kj
���:D:5�SF>DM�/��R	�t�^����ZyMл7�C���/KM`��h���qY��M��S�o5҄�{j�
�/��v��>�P�7��| ��wVE�6=E�$�p{��svr�\-E���x�zX��\����C9=�h:�zs���78����԰��p[/�y��\4W;{���Er=�K���+�Ɗ�w{O��� �,vIzr�u��O��5Npj.nu���,i�����KQ|K#y�����Fe�� )�A��♙���01�٫�z�7�4��-�춡��w�SO1�Q�ul8�G����5�$� �z5��6���R�����-��+�<�=(�0�1F�yo8
�\�&/�N���K�v ��cs�Q�:���'�ő*%nZ�b�`f0G}��76�n���l�F�#�D�� [;H��.a��=h����hH��6(Gk}��79�~����S�2e���
ǯԏ�^�~0�
xD-L:*��oݛQ[��ohW� �l�>>��3����-eCk��(琥�"�5�	�\>����s
�~_��-C)�s�P3FE����M
��9>�ڏ�ݪ����*Q�ӜH@)x�X�N�U�u����4�Y|$_` ~Y�l��c]�ĺ\��`�+nQ*���eEK�PP�H�Uq��Ei�|��������ߋM�uC�_?�ؖШ�ִw���ؾ����^�w�pz�A�
��OV(8�̷}R����G�T�Q���p#s�w�iKB{i*�	(����"�&�u��V��#з����>��;J�c쒧��5 T�^8:xƾ-�|�"��i����+�b&Йp
��\�,fYW i�
�e��5��8����ʙ�{��@:���A�l@B�B\L-����AZ�-�>�I�p8�>�;5R#^��_��`���BzϿ]tzE*�b
-L�_����Cּϔ �4.2p�vr�r�W��m�	H:Ee��x��^�h�c���싀:���"_��;��TTsv���S�T�z���K!+��7�$���ߏBO�D�*����c���L�=�gy�J�v�B������Lo��������%��hav���������OQ~�Х7�kN�y�h�ߒX�1�1bQ���z���s��ɶ���#n@�f�i
���//o:2�����q�]�1#�O���s��$���GG�1z_���ʱ9���-��G�r��q]��b6Ü{/�l>�@ /7�.�D_v=�#XI_�H�����5;�kR���G�����5�	�P��:/|��5*���>�����Q΂s����8�ܑ�Al��V���<�==�X[rAYƫw��ė�7v{4���٬�U|ҩL��p�FV�>}�,%ק8����itB�o0���� ��+�N�E�;=��9	p�p`���񙐲b'e��L�06W5�w���MQ&D?3��Ty��N?�O.�ޕ������:�Z��~1��*A0{ז/UR�԰����A��CU ���
�E׏�D1�h�`VY'9���Qp�cg��ȃ��H�āe����:�I�9f�/��xJQ�cJ���@r&R�lG'�ǉ"�|~� c?�:7������P�7�.��W�=���_*l7�sH�]��d4����d��r~F%?��yկiwߒ]t �dq�8zש��l�v_#���(�C�����ٮ��',���]3�a0�P�l&���X�i�`vu\S:s��e�N�G�h���� `�9 ��x�r��3h�����܏m�#"}߯ky��BH�����!�2~鑡�j1�F-�LG*v8>օ;��b��#�wet�"�G��b1>u�s����ᖤ�_Q#ɑ� ^��e�C
��,x�g�w'�0N���3���5:�:�^AF�K�&'�h��I��h�,��\�f�:y�V&-�^�Ϣ�nU< x�[ӟ~��˗����%V�b~Jd~����9����6�IȒ�ѕ"��(
�t� Auċ�.�?i�@����[t��^��c!��-	ǫL�yJ9�7^l�''�F{���+9�k�y���0����甃�YRt��t��@~�m���������T��u`�뎯v����p
~��g�ު��� �e~�GQl�����1�Oy�΃�]f�R��ʂ��e*��غt5��l&�)Ȥ"��q�=<����*��
�O����KiS|���׊;�����0-��	z�O����u3vU�Ӕ�� ��|��C��������*����J�Bb�d��U�&#J*΋�̀[t:6�ƫ`�2�=��-4�hHd�"܋F���ۇ�J'�9��