XlxV38EB    208a     6fa�A�-�xW��� |rOl/�	�u'9��� Cl٤���|\�(��"/h#!��ǖͪFw��8�UBa��p��S�,���7������U�����(�����r���|/�(����r�i�_w1R'��	�p��r�vm�CYp��グwQ.��"F���6���^� �.ΌB3=�c��'�n���Ǩ��]�J�Vk�[�I~/ؔ�p2.�g�.��_�r�6��[y�� \�e��޳�(fE����Rَ��_�u�ۧpm�v��8C�p�70�{陹	��ya*�n�a�fjd:��J߸�ԣ��W�KgT��&��>�s8ߴ�P�p�\3#{j�䂔�ۅœ��7f+ժ`�Fl*��A�)# S��d�c1�����d�cV�=�رT�!rґ!�p�nێ�}�H�Z��PI�j?/Aa����V�hA��Y2*b�oUL+�X���"�����H4d�jf�	CUr��N#���������\��ox	\;��4�('_=;��g� �z�bZ�f���鍕������}nhfu��UռТ�N݄�OE^l�>ʍi��di��<;<���49��x�/1y�����Gu�1a(w#s���7��5߰�������O����L�<���v�z��Kg�m3F�����Ur�+�}�!��7��݁������hK�Ee>�T�u|.j5�_�y� q+˧��U��Y��y�!NUNӖQ>0K�h鸙��n��Fd��-���SW��_	M���I$��^QƧ�Vg@mb7��]4
�S�U�H�p�b��%ål��)��J���aB/���揖�U�ۯ���%��S-˟���>�-�;{W�� F~��Cl�t�<�`�T��j[���+˛��k|��^G��<OV_&`�,��+��E�2@]?�-,)kZ��\�M�ʎ��4�,ǟD�����A�,��[F�r,u�&|�d]:Q�0>�u^^ԓ{�kfۭK)�HT��V��m�:v�x��fX����9�z��E8Q�x�vE���f��~�F�h紿A��E{m����F t~}���t�"��fy+/�7�'zq�����Wn�>-41�!.��6�}�@\Jf"oL�0L��Ջ�.�e��lS=/����l��FI� Y-���ٜ��g��� �E�X|x�$�e�s�/1X�
�ޏN8�Ç��0JW�k�+��������'��<ʒ���̦�J\ O�6���Z�F�F#��lO4�F�̷��ZOlH �䘟�����j�|`�mTR}|�>���~9������?m��87�D����$���U>�����u��/�*m��+2.���B�@��!w���O��?\�{�c�uX��{�à�������Y��2eJ�j'[ioi��A�G��'�	'!N�����$6W E8�{P<P���-B�o�����B�L��Ln���[���JK�2�v�Be�_Y�8k�#�T���G��������a.���E|�&3JdŖ8~
�Ry�A�#�g�:��c�#K?�^Y�:2�� 򙈦��-���L�kn	ӗ!ݔ7Y{_� "0�6;
Ga�3�퀉�@���?�:�t�o�oNtc�{
�f.7B`=$�d�jzDՕv��Տ��
�_k��E�����5�6�ٗ:�)lyq����?����I�2Z�uT�/a���� ����I�י�<{	@h�{o��~`�t�P��;ܷd�!�w���A�LZ�}r�l