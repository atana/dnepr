XlxV38EB    3a46     8c4n�."Q{���@�NרT�D7	�Q=")���F�&�+�]՘B�%�; `�X�\#����n��<��Eӧ��dD�sg�|Z����Ƃ+)		�Ľ|�k�L&iI8&d�DWQ�@ʑ�з�@�	�J߂ML�W�L\��Ϗ�1�\-���s+9�}�� o��ޠ����C��'3����X�+U�5\�a\�����mm�RP��f� ~	iJ+��Й9�P����g���3f�b�I>�i-���k4v���<�m�J����{dTr���8"�� WGΡKpTY+7
���Lw*��-�C(f��~U���Jدi���YI�����t�V�J�䬱@����3��T�V�K<�=˚*��)u�a�0�jrZ�߹э���<J�8��ad����XX@#�#ۥ�&A;Z�����l�{8s�J�Yn~�SդE|��(��v��i�����;L�a|k��I�s���[Z ���_�#��W�"'�'����R��ԏ�S�&��ƾc̰}ԃ���Z��[;�\�m��w�`��D�NofR���%�(�v� ��ں��WP���_�ʹ�f���(,�(�#�d|4.�Z�+�2aL�0ue�Kk[����C���1�p����b�Mg�C&��ȩY��qV�t��_����(k]o�~k�򟮁c�hx9ƅ�����)(8�Jע�̟��KH���H/�ȡ�c�p�{��C�;������J�RI��q�a�l�(-R�fN
@j�h�U���֒���t_E֏�]mc�p.>�%/�B�8q;�>�}x�Ј��mɛ�1���g���u��r�!�Òt� �,,�u�s奋��d�4ʹ��\�a����.���k?A@��U��0�s󘶴`�x%�_��v�S��-�_i%���+�g�P*��w$������}X�ls[;|t1Y�Ŏ:OB�(��G%�8�龪��#?��n��4���b���C4����9�)��u�樓kBf��(uY�v=l�6��p	s��`������jc�jt&����Y��Qjq�L���X��2�t�@>�6~!���b��}YѤ�v�qt}���%n�
��2st�]3��woa��)5ji�du��Rt�����<f'^pUg�Cr�Y!'��������j�]����X��,w�Cau����q{����T$�ׁ0���V�4�� ����w��bZY��ۋ���/��[�A߶�,���H����(f���a�N �Lp�¹���)K�)��
SX�?�ܿ�ܐ%�)Y	�g\ �+�zI;���ϱ��ӀA���A��O�s�rX�0nlB����Ӻ���oc���6��#������|G�c����{*v����1�:e�qW�
vh޲]5�P�5��VK�}#i�܀��[��q��蕽&�R��+^�C��Qڿ+<�+�
�W<1@�&F�
��M3�WW�<��TV�?�0%��
�b�<ȧ"[8�AN.s�z�ݔߨ�,�Ᏸ@�0@t1e�+w˩jE�ٌ�#5�pf�xp�T�Dr�����D���yd~_!g������k5�v�晳�H`(�����ثq��&������qa�J��$�=�T�@��D@{j��ӿC7���!��6�����$RRQz��W�<}���dɛ!Ҵ����&}>�$�7��!G�q�
Ѓ���Iby�=tsI��(�8�Q�*�N ����6
�.��5�\���S �(�0/y(��%kƨ����Ίsfva�(�	�+���ܲ�IZr�C�ܳw�kB���ޣ�>R'h�TM{�� ��MSNZ�/z��O"D�؞��RyWrEl+N�W�w����f��=�1��o֣��e@� �b���Z���&�]������*���ܟr������l�#*8m.U��O�~`1�(�ϙ��0�흝n��S&gtJ��?���]B5z��f	��F4{4�H ���)�M-�2�4�@1nT����5-�0��D�n�`�ypl�"	 l���
ߋz��Ҿ����N�c�cx�eM�J�%�
T&��s�8�A���*��/ڰ�%�V����:-��G��ڋ#(�ڻ'��]&RhF!���#3j�Q]*��Xϗ��s2�%^z��@m�.|�2S�]Z\3�v��yU5��y�����X����jh7P�0��[�������O��D���/��,a�˒�ty���3" �zTSB�