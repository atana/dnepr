XlxV38EB    23de     74b��6Ϛ.P���K�ρ��l��ؙ��Ħ�p�KY���J�Kń.㰊b���)���_E�v�RF6o`��[;��]f;�6�������k�_���;U��-Z�F����>���RΓ���ayt b/O����ƞ���ٙ�^>�k&�;4���Z���)��-�R�7���N�N��雽n(Zr	lL�����HVo��W��}��;6�Y���w� ����N�)�<�W�+��	����"�y���c�-�6�֫����c?��#~�&�T���ɫ�i��syJ��A3���g8�$��bőֆ�X�_�HEZ��SÝA�ȦŹ���~L�4x�ꁋ�.� <�a��5f�.Գn ��
w��c#�[kz{�=*�HK�>�aP� w����ES^��´k�.xNWc�[����<�k���p�<�MiGs2Z����F��i����W����~=�O��X\�X��K�C�+q��b�ɗGQ�v� O�H]~�g�����ݤ��������]Y1�3rάˮ?�R�^������s�s�@KǺi�<��	����e $�ʊ�K}��U��2hl�gw�e��(�����8��x�X��N|��4����]����7_b<G]�ü���Qr���'�X�	�����D�2N��"#	�`��%ȑ 9�x���l�A�կy/��V���g�>���h�uU�W�,��.������ಌ��␺�׊��\D�y6��$�N9>�A�k8���Y����ڕN��b���WA�g>yFtt�c���~(�E���HX�/��+Y�� q�c�$E�+p��/��y��0U.�U�MY'm$_L��2���[#��Ի�<�%ĝ�z�_j�#U��ê�����`�m�6�$E�73�RSy8"m��~ui�ωM�c�S-�]_wD���4��������,t&�"i塧�C���j$X��Ѯ7�W�)ٸC��Ux{i�J�A%a�m�Wc������}-E8k �V����跴��� �bp�p������ʃ�D�@lSWh��)n��]�*�Ķ�(�9h3�[�x]k)s�xYGɨ��i�/�{��_��n�ũ�X�o����U*����#mJL���^vF�����ؿԝ��⢿�.m�@�~ 3'[f���.7��Z�9ٰcو��Cf�SޣR�H�U�%��`�S.v��Y0c�[S�)a
yOtB *$l+;\��fjfFĝ�f#ƿ~H8���T�����. J�PEO&ľ#��/9�22�&*ad�$l�Df/:�XFԴȚ�(��P=��,6t\8+���N�\V�&������O���M_b(�6��3��~�P����,(�f��,�����_�Y��8N�E���,���I�R���t0%.~�-@���5)9�T�����UG�ۯP�k���w5�N:�K�{)IM�ݱ1�a�S�9�>�پ��=�2�W ���ƩI�����4�E-��K���텳}G3�cz����8{��`��
�h���VBqC\��00�4�0*(�؀ڻbمN��3 �L�2�P�q��;
cP�آ-G�J9u�s�Jg��%�6����ěl;����`��1�S8��u��m	���2��g� �@���{��MƆ:����˄��3���	���ã�?��zz�`�ё��'t��8H���+��%��n]�lI��/���lX�4��vh��k
��-��B5	�
�d)�('��>��Z����Hon-%�G�bƽL��ƚ��j4.w�*�&�b]���Z�L;n�5�\�A7_iJS�P=v2pemh/�\a�n��Q���8<����|a$^a����H�