XlxV38EB    10f9     468�пx�k车�5�P�Qz_�d���UI�%��������(}X1T)Cll�$h.��k�f�n���f�	� uk�Y�F2�c!�&��H��$#���fA		(��d�9�t��&;G:��㗗�3o`y=.��2�{Pw)�Z���pJ�}�v'9�}��E������1-�+YږJ�&@��.8A��;;X�85�;�n4�p���]opo��O�Ym�@ZQ����i���x_{���2�=���8=��6���#��	nkh�R�X�oDX�g���?�bi�G�����T�'U���2��� �d��}m]1x��>��Ч�,�'��Yq r���3�Iic�DxM� �K�T$|U>P���,��p}�t`�ĵ(���\�KQzB0��ד���?R@���N�M|1�ݹ��ZX����fĉ0�kc�8��I��CPI �������� [�� � �#�b�Rv$lk�"��|�	(~}�si
Yu�b�~���3�J�$g�y=�zzko�3\��4�f���qs�� ��>������"/�����h�4dT��ЋHg�4TV|���`�W�)�[�i�9Qႀ�sz �3{ԉ5'O��)3�d1{��	O�l�g;g�ʟR�D͞}�mC��ۑ[�'W���m!ԫף�<��ג2v�"7c�D�WA�9���v�Y�>.�5�Z?9`���T���J�:�'<XFVȥ��?)�E�Lg��9$p�E`�A����וs�պ��pB�h�����#ǑG|q��cV�~c%z�uUZ�A_�et���p�b�P�|��Rt�u���ʨ��x����9%T�\6�v����}�vR�v�\	_�G(�{����5k�xq���&(F9ԭ�d��m�Ћx���Od٘[�w��$9}r#0%���d���r'u�:��q~��	]�ajLD&�F�HK]��瑔�_��|�6nd8�l82��_(��>Nh����u?`-��3J-k��%��w��5�~�P����mm�Ա7��[N��*�Vb\K��o����ѝL(��~�SM��9<!+{��4��I��@�Sx ��Z�M:�֦���Է��������=1��w�����M����^��˖g�C