XlxV38EB    8d4c    14c3%�p�z��ii+�2�.تt�ÚRw�P��˙���Y�|p��qN#�&���C�V��D�DG~3�ο��Ň�!�.BP�+Q�~�E���o��r��n�UoR]���e�t� Ev����M� �����%���=29��.��mei�g���?
2rN�\N#�"�e�����|/���I]:��S�	��ǡm&�d�f<��sCϝ&l�
��ӯM�"$d=kڠ�x^~J�J"�7x�@s��t�GQ��C[:V���	u	�Y�N����f��Ҕw'���EV�~�j�4PH�R�捪Ҍc*�+�y��7�jC��nB��<ܕ��wꂘz�B��Qe;9��-,n�Y�t�A�@Il���A�u4u4� ��\7K�b����j��&��"'��|ǉyvID��7�4��^%�֢���V�`F�0���1(ID�0��ӽf<K�
4�����ɝO�4v�L�j.�_��!�Z��a=�H�B�cܞ�9�bh��;Kxg1�qsm����%9��[�J��@���q�>��ۂ�5�e�J�=����h�U/�A�'p����d�������X��2���Ҡ:�0t݋@��44�tn;�J�>*���%d���۲�S:�:e���]b������
 UY���E�|�7���:}� z�i�M.��7I��nK�Y^�� �|~�4C�uJve�N���3
�%�aH^�kx�U����ۍ��.�X�G�=�|&$�g;$
�yW����J��f�y9�)���/�������׶!�Ə�&�q0�57B����j(�p��:�[�7#��lܟ�O+���ʯ�j���.	�c�o�l��u��W�s�c�S*+��D�yi���f���~��&�
g⌵�Ŵ����M�/Ĳ�2H�����$�2vv�CNq�p�X�P���6��k�dF��[�U
&طY�%��Ș�ҕ٪k��LWRwFg ���E���6�Hԣ^�"������ڝ���B7R��Q�I�f����K|iL+W�V����Z;Ǭ�fCy@|	1��[���[F��������k��N�ґ����iǅ7���2��B���`��c��9���p~����7���@Wn�O=�j=Jԩ2bs%���%b�� ��(C��Ve��p�	[�����q�:���Q��oMTT�/��G��{���B�E=��_q��{\�m��Ŏ8�X�g�>J	L�J��ᅚ螑�6�Il�M�:��h�g�׆�i-�NL��S��Z���j<��)KT������(�����3 #�"0ч�@z~�Do�-l�=��(����
�d'wIo3����"��=��uO��PҘ����hL��l�M1��~��13+-[kV�d?���ԇ��+RJ�ID�D���:�	�rh��C�y�^�$;�~�s�Z��Xf�䣣U��VZ7�j\Z�_�ަ�R�M��u���^<4ў(��0�/A���S����(�m��<)���A��1��]��J�9�bA|�]-/a5x�H�n���{w�����i��d>��ea�S�>Q�,������a����e�Y	�"#94z2����a_��\�ֹ �
6C^�#�&�B�I��v�"��F��^��օd)[�r�W@�
y��w=^��l�����*�D��o`���W�͌xT�7�[��ȟ񷨈�q�:���I�6��;5u�í]E�YPE\��+_�Cp����R���G,̓V��ݡc�<����2ե�������z�9�$ULpU�3�|��b���r,Y	�����OZ�-��w�p�Eݳ ���*	�ݐ %�YYS�[�ւH�����M�ݞ�fL��+1�;QGz(D���E��������u2�itn���5�d��)�*�cw�Wm��:�w��g|>��Y �Y���탮Ǹ[��{��6���:S�	��0y��#���ل������?�E��1���n+�,Wυ[��ͺ�(T�nD>�]�V�u����2��y�7������
@|at���4��SgcP?P���A��C���Ki�Z�Dv�B���TI9�=��C���r�+#Ĕ�#Ғ6�<�9-�[|h�K��<��H�!��3�a���?0�x�̴����݀�s��9�]|��ee"����~NF���}��`�����ThVܕp"���D$����{�Z��j��U�~�C����~B��XԸ���z��5�J
����z'���@|/�R��u
�e�1w�]!�_��O�����S�٪j-����I������R�d2T�T��t�h�d+�V�^?)�����wc� r�ſQl�!8�"ÐHe��]c8��xB�hgw�A�^۸9+ʗ�p��ڀ�c� v�����X*�3�{��|o3�*ÓJ��/��{+�Z�@��Q��,����X�d����|�w۔��Ƒ�?K�år��V�Ⓤ�V$�(�ݟ��� S%�|��p�����m(?u_9/Ko<���Z�X�d������*���8i�G��u��aLb����%��_ebq��3�!7h�<�[��Y�Ppw��#YS	�\GJEX�kyI�;�&U,��,�W�9j���g{I�[�!ʢh��V�}�^@�L�`R���,����$,��r�%���)�S��C������ոF&~jE]\�r��G|r��׋�^��vOC��rs��Q!�rk��W/�[oaU�5Ki�Z�[�x�qa+n��ד�LϹ`�`MHM���4��n\Xar��:O����-*#���Z�\��-A^3#z�ϥ��@r�7�چg���������Y����Ʃ�B%R�����&�I+6�l�>]���Py����Ļ�{ѻ��y(�i+�����ݚ/YG�{�~�2z���Pu�%Szy�[�2�������d�x��ۥ2��Vl��-����&��i�!��qn�Ҏl��O�q����hc@��,����mQ7�m�40t��W@�:R��M���T���ixR��oO��N�#��� �����Ä���O���<��3�<��uɘ{z�w��Y5�:���fu�(��y�T������\$�?� ����_�Ʀh�xX��/�f���c�U�x��/������p\����`�K��-Qi�����ȚS?#���nS�aJ"9bTv��ڟ�[�2�"+���kD	�so�����T�!�cZ(K��];�K�TF� �,.��gzUO۫��"�|��X�}���j<W9�����V��y�xǊŴ&�/uW^��� ����m�os-]HHUVb�WS��)�S��M��3��w�\�y�����zz��.,m����X�^�E��:U��}3�$��[���PZ~���p��R��z�	��7�ԀHd����]��NY�� �];����F�c��6�-�>( �p�i��i��k�����Zi�9i�Ӝ��ιx���M2�V(��,*`2��� q�K��v!+�͖ݸ:����E��3�5�=��`�U���z��誷��Г�f3Ҧ~?�d�]r�M�#��GH/�|L��S�����ԁ�N
�����*�C����&����iH�j�4��S���PPm�A	�X�~�����NZp+:��y�ׇ���b#J���2�M��YX �\�(�6d����diЊ�3OV`#W�D�W�~!9�-y&��6�o�2'�cp���_W�� �����Z����?��c�r4p�C���d�-fu�Wm�o4(����$�LV��R����ub܃\K�0�?�txL� i���nވ$7@^������4��0@���Z�5tݞ��D(������ֶ-�/iwH8?�����zRG+�O��{T.ni��G�	y�v<^Nע�PSL�85NY��n��1�T=_��)��A	�k��liGǝ��>J��vꗮ�=WxsB��X{1Y��4׉��A)4:����<��wS�h�Q$��%ݱ>E,�#�g-����+я���tRh�#�m�a�q	��@Ɋo��&��?���c4�����-�`��j@HE��E�-�CF��I(a���B��~�_���d!�}�mۀ�wdg�h-4�j�z��X���T���vK��:����ݷ�����b�Uhx�!�ݒ�~Ug�����9��Caa��g�@���1���E���O]�c
�$�5�GS4?;��H	괛@����J$�>��F����v[�Y]��	�Gu�hS�9H��U)$�
��8f�9ۋ���*�NET%5��R��B�0�w�Oѫ��6�3/�O�R|(��?8��ڥ�&��'��_�����(L��S����К��D�ƈ'��(�����-�l{5zy^x�������^�4�̹�mD$�4S��NKl�v��oBI���c^�%"qf�~� ���	�P��" ��J&��j5
��G����F!�'����� �W�r8�(�?�	8dNqU�Q�|�nJ�����8��/l�^tV�ZL�y_�G��m�������B}����G��IV�܊$ G�s�J���0���x�U;(���Q=���o��I�~�evbBsUӜ8�V���Gt(`Di�ը"<pi��ЬҲZ��2�8����ׅU�:o�h�~	+�Kߍ�p��H�N����6N}Z(h��GR�u!�{E?��.�F�xꗻ���@s�� x�=,�gD����@�2�%��iW*��tKF8�Rݜ���hk�e)�/9�Ј���L�N�	����[�0��)=2��&��{cY:��>����U\�̐z���p7%Ur������n2<^�.�G�b��{�,�Ş�߫g�g0;�����1����Moq2��ٖ��������X���,�#>�R�KqM5'T��r}i�(Twb������=�3��[lN���|�$�J����:_�������_�]��頧��i͊*�{��� q	u�;�����6%���+}�M��:��ˀ����IO?ϗ���`6Wi��f'�+Vb: ��k���x��3���?��'rR�7-L"���~�t�Y�Sl����3�\ʥ냓Ù���AkPύ�B���.��q�%�z5���,75jH�Y�2�*��e�݌67U�1s)DXKEm3k���{.*}$����G8(w�k1�i�C�]'K�q��pM��͐.�ѹ>(s|���=q{����6r8S�6�� ����x@	���o�g