XlxV38EB    9e1d    18380(�1�7�&�*y{���S�S�ɚ��Uj��:7�b	1�{9����,��xp��u���@BJ�D|c%-��B�i�$^�c���6�ٴ�
 .�� �@Y�XX��'��Q�O�oD��n�4҉; �yo�b�g�?ǳ�˷.;�,�� ��7s��8��u���'_{)N�a��ȶ��3i�p�$!��;)�+�Dm�m�}1��u�ڽ��f��f���쓎5��.��d$-7�9�=���|��v�1lhY{�*�1��u��DoQA���U���&��;?1i��ᝌ�d�F��d���n:�U/�Sĵ�@JM5����t>4���-�K/��}Va�Z�M���I�0O#�h�Ÿ�3�Bb9��WE�k�{��t��<_���(�mu�y��o�
�Y�Բ% ����	9��ݛ���M��(2;����ʹ�n�:O%i�ZnC���vU��WU��`7�٦lA[B�G�)k2�̶�M��)�$�I� G(ߍ��!l-�QЗL��"�dy��x��}{A���	msj�t�V�y&����(b oׄ剠��#�+S�{p���=�d�x{B�A0�2��m:����x��"	����\��D&�P�00x�6�s ���<;�����;��B9�䲩ظ�.M*;��֞�'��-�D�˕�����]�{��=���'���nG�'��}���� ����f�ja�oNYE�s^��^��2앎��e��:�}3��PX���6f�ݻEc��}��]�\4|��g
&r]hZjȻ{S�CS_TJӬ9��x�F&��A� �*��[����2,�O6q)?;X�����U�����N(򵛌 :�:�������ٮ&��bW��%�����J��S����7}�t�I=!n)���"�NG�O�y(��C�)�`�f��U~VoW�3Jx�LZ���XU�7բJ��06�,&Ҭ��됥TY[/�K��.i��׷+d ��B�X�J"X�:t���O}/Cڀ�<mdu��!.ށ��`�?}��b�G'%p�|�H�JlL������9�$�l��";�ƞಧ���<
	�*/B�w ���;�F�Ey��#�P<y��#]!E�e��ahyaE>3&�<���)��f�ؕ��x�o�a�x�+���!Q�����E��͒=�EW�T �!L�m��2�ѯ:��nc��W��52;���_�uL`!�C�}�� ��H�W,)��h�3��V���4b���j�[��I)DQ,��Ƣ�4��nf%w�Ǽ�>�^V6)���`�w�%�{��Ao����� �ܪL�!��n?\F�D?�-�2�(4�M[(����C����~��c}|���q��a�)�-���͝�	�W���/��F���m�-$h�;.�-;h!�J.5�̃K`��H%��<�[��+S_���g�����0�o�~�2����_0�g�	@�蝼��-a�OX?���ݒ��m!�&��``�i��96�v�X���)�˫���|� A2b�;�t6�߰�o��B6���dW���ճ��>����5����l�*��g�zǧ���=���\7h1:���C1d�ڗ�:/���Wn0\�D1_�p+�)���g�8�����Tj��F������5*�F0��r�&󕁒�q�Lk���"�O�������ЂF�7���?�ݠ��UY ɩ>�+��� Ե�4�Y�6�(b?��<Z���2S�<�̃�hm�a�Q�kU�Uꜰ����;�5#�5�������}�r��z!��Jl�Ng	Rt��f+�@>[�-e�C�f���ƹA7LO�������Ƃ�J(�C�A�� �853� o�>��2��u�%,�{z�N��{��!�0~@4E�14m[��A��V��^TZ�5:u�hV��uμr�py�ʛ�o�%�`�/a]!f3��(-�װ��央Na��c��(��̓,5W���b	Ŏ���ênMv��彋�&3�r"K�bZ��қ�8(�i>e�"����r/��j�u6�(:���3�i��jю֠��~�ɏš�J�hvB��O��f"lͪvI��3l.��&�~�Ɔ@4���Hpq�E�{��nҔg�ܖ���L�&�]{@��5QB���~��I}�n��Iz�_tS����^ex�}���GZ����OV�n׫�� y�Ƃ�Lࣳ����i��b7�_��ӿ7�ê����g`?�I��		�6�w���zT���j@th�A 昛�y��W���6��u�GV�M����('�F��{��2qTK���ّ�|lc@zy�D�C�>��O�q�����'�X���8��1�c�K��7v9;��}6��:j�+�攙%y�8�	�~��ly#��_��y�O���M� %+C� ����a}��t�0/����Ă!*5s��R�_I��Н$_� ��]�Y/W�7v^`=�^Vr�M2�Eա-�x��GK���Q��?�����!���p$��������8Mx����E��s���WnK[��^�9P�4GxE��� �<��Y_,�޴(%�0T�A��	٥��`�l�������
���*d��p��(�"b�"N5����~<���mܶi�1����)���2���
��B�p���_������f�A�����K�2���t.�P"k@��{�S��"���K�2:�3�7d�k}Ϳ>��}���/�>K`r���s��<��d˥ӑ'���-��9<�`�d3���"GV/�pײUӗq��x�����@p`Y�q`&3ʽ��;�_=�@�by}�z������F&��)��|������տ+L=j.G�.:���<s�T:ߘP���|��[}4S3�/�f	�&Ŷ��<�%�J&NG���޵qʼn�F����n�V�"�#ǣ>���Vs�S�	����*]���Z>ںu��>�s�*���Lk�/��ќ���;�Щű1�縜1�M�!�1{2��3�����N�.���x��K'� �&����{��	~1�Ţr�f�ͩm1!�9�ݳJ�m/cwnK[.�n�5�Y��ݪ�'�qݩ�Cw.�^]��y0��v@G���;��>	t�Ga>��������7��$����\��G��d�4�5,]	��� �{p.`FF�=Z!��}�h�1���㭛���'��U㴣+�ip1o�j�X近��D�+����r��?�$*�<�umM�� ��K�X���c�Ze����&����FQ�|QM���R[�t�G�LI
�>Y���A�ϳ����@�5�����F_�7��d$P�f�:�bF_�7��qCv)��*Fz��27y���ԓG��@�%�c�S�9��KJPU��BUߪ��[hL�c���1�u���8=�a���*q�TŚ��,��2@���a�T��@��ߎ���D�'��}�C>���Dsa�F�~Q)��R����v��"�F��m��N�m6h���������B���;�y�Oҕ��5�j˅�!�F�`��7|�|�-�'�у<-|�M�i�+r����3�nG֔0�m�=�oe�0�[Gg҇�fxzX��Z�+�ۅ��忊��������ڰ�s?�A:�
N�-��'�H_�y���oS��SL��x|�����-��e�'ǉ��S|N��޸�
�R��8�J��L�[��X�-��-$5P���H���� /ȥ.p>�pJ,k�8�.��MJ=��l�y&��׾W>�Y�Ѧ,������[́B�d�.�ॽ��"�]8V���8_�J�(%��4Ef��N���D��,iH���<�5@�V��6����ɄW޽mM59���P�]�A����&H��C'A���c��/����囧��C��� -�tDѥS�)6pa�9-���m�� �4t�&T�J��n`Ѡ+�����6`Y�"*=��~���徝�64���o��ֆ�rq��9�'�K��Id�ɺ{�v�1���3�w�4�����s�xϥ@����<xIM� �L�S��%e����Go���Av������L����&4�~ϧ�3X��E���c�m-��_������]0t�3'G��N��Rw[�����}�v������I~GT�+����}0��d���Ѳ/�j���;��0'����g7��ӫK�%6���#uh��n�j�g5\�=���V����&��1Fmj�ŭ�Ki�9�ڦ]�:��w�
Ɯ�풷��ɦí*�V`.2i|;1L�S�h��ak�x�����'ņns���i���U�zPO��1eN�V��|��=��6��(UHV
��*��j�d~p-����&��uj$s��x��iF��r6��#��F@��_5n:T��~�N���k�������\l�?�'�ȑtO���s�y����
&h��b74.�a�����;�����z���؅����W�W�j�ׄGd���k�mzcS��0'͂R%�.�����|k�S�a���p�;Y��`�u»�;T뿹�Y��C�_J�\MLi�{��Bn�;�6��wD������!��~V?���b;�����^..��~�Z�W���Yvy�0rEuo)��6�+�;��۶���e8�2�����9���h��S���jRφqOG%�_a9�_��8T��P��m|
�j�L�4Q��(ڣ��pׁ:��#�SY; �{��*�ghX�M���~{>׉挹Uf���U_"�4%qMu,I��4y7�e�d�Y@D5�p
�<B�˭_|{AOAO3��R$��Q��~���"Z�����ɱM>��ܣ(��?D���,�l\Lś��-8O�2���*_O���f�糆��x�7W6��P=?�Cr=�)B-ѸO%cgc�Ak��S<7UΊ�{�'���-114�)g��K�p�#�:���L���1�M�Cf\C�$.m3o^4�ۣqؽݺO�Da"�3G���P��h��b:�o�1W�;@-�7`;R?/+�(J�R��	26�SU��b�!qj��21��h-��w:��8է�rU��}��C�v�O��ю>}�wN��h��Ŭ?�L�4���D���<,��A����5�?o��]��U�f�w�$���3��~���[(r2�wM����w5��ζ@�N�h�2����/�֥�>�xׯ_k~��v�~����{@xA��e!����YC���? ���-���C���/�Cd���@�=�	b��!a-���g"$����aI$Z��@z�o��2d�')��1F��1��Ȉ�����%N��5�#'���� 3M�-Ҷ�[d'˹9ݥ[���:o�Y�?-QcAk���`v5_Us��:[�O ��²�CgSn�3*y���H����k���v9�Y
��8l��b"(Z��d���E��9yO�q��,�8����l����ԾzT H�#S�r�~�~B�"��k  ?E�x*+N�G*�$J�Ѯ>��_;k��m����j9��m�?½P��<p�� �}!�Š���v��8;�n���N����on����]�t$aQ���Z����qb(��� HIO�$��FKy�<_Zd�jW���3����TȚv��Q'��D&8wJ� S�{~m�Ql��Qo*�R���%�es�g����g�A���0 �Z//2��CB9�6&aѭ��4?i[�����F�5�i.��"���}w`�a��Ð��\b��\��WƆ:_�ģ�]�P*�k.����700H��$��W�T�xL��_,\��M�C��R�Wתd-YWt�����7j(ޱ|
��fJ%�$Q���(
J����䩽�m0[~����
�L�n�X�]����!c�Ma>�������I,d�=|���*���U3���
�:�B�Gf[{w J�%w�>Ҧ�G|�}I9'�_�_3z���lyg�����/�A�#�����d�\�=��4����:&����=@�W�]�c��Z���^�,��ϷaY��B>�?���&w��/.ô�;��'k�dPA�/��D���z������6E�r ]�[K?�5 �l jr��3�.�vFi�|B���x�:{a`�������\qn��$������3��'�