XlxV38EB    316a     99aUxm<Kܶv_d���"�(�E�J�K��ps�	��fH�P��uV��t���������ڱ�t�t������6Tpd^~�D��yX(��%l�T	r��`$����"�2�yȍ@�Wb��3zN��l��Ie��Ԥo�~�8���=c�d(��.ZtI&!�y�+��2��\��,��Դ[��5�*L������G��K�{�S&p�GJ��j��:�aDS���J�W�������H.z���R>��ZK`=N2�0��+S��ghڌ@�<�������M�dK���,2�l}�ʪ+VqJgG�	�J3�o8��*@����r`��_��	�,���k�9Qf5w	����Co=ڴ��v#�_����s�m�y�,�����#��v�Mom�d�c<r?�dt���l����p�a*ɋp�La<�Ղ=��,�;�K��,�/�-[�I��;�l3��Д�K����\;�h��^���t���b�B��s�P���=��kI�j�#x���B7�^���f���߮��dЉ0j���r󕋍W��b�7V<�g{6���x�|w���.�+�H����-H�
�\����k}Uc�]1%.p.]���.��djOM_��=��ڱ�Fpl]6!*� ��8���u�������,F\�5��(W��HW%����M����>=x�y��4�ؖ@�;c9tn�㎺t��0�mk��N-��&p˚����?\(	@���=����p</D�2����s��(�pS�U#� !uiߛ��-��������Ȕ��w�YyqOλ~h��-2�ѕG��u�\SO�,yR�j���<�-K��@I��>�+N$����^��o3�A�KF�f� ]2֖7�T{VA�>���븍�l��Q����H�h�9�e���c�����b
]+(��x��O΃%���з�S'���� &O�C99�I��¶^�N��$Q��	��&�%8�Nnzi��X3��6�7��&�m��|u��G�w��8���sw��r�� eR(���y!�Ř� ��3q;*A�xߛ~��z8�cO���La[Bcl,n�/���ɪ�5>�P��\w�w #RP	{	{���T��*/��o�|�w9U��L�\'M�`]SI9�Жma���b�N!�����/�3P������C��i?�K[�.7 �T^��x��00��3\T<��C���m۹C#�
��Z�`��;?]
'K�Ň$��?c�*Q��%�0��]Qk�I��r�3�Y�F�n�1�5�"��)��=��n�c=?c�Nco���Yx�v���|l���j���\U:Ŀ�ݠ�fo����W���T/�և�FV�<�
@t���ho��6G����Tc��r7��Q�һi�|曩�[A��I��m�ǽ���ʭ8�
ASKΝy0�l7H8��s9��^}Ʈ���"Z����;l$^��b���x�I���B9_�'X}��JHǡxe�4D)Oť�Śriܥp�1���������:;a�f�&��
�O0�} �Lj�r���V5�,DI}{l���.��� ڹ�"��1�IGtr�����c�k�w�".?�
�A����FuuW��²;;��o7_
���[c�έ� j� D�+ApO�JX+N.pasD��8&�؁In��C�π�����g�C��M��xk������_�aG���V[�j�h�ޚi�������4��Y������B7%��/�$SE6�_)�逈Bl�T��I+�w�Ⳉ�>�Es�gh�!��T#B����`��(��t;ӥ�?2)ˣ���ghM��zcZ��w�kV`bg�
f��s�L=A(����|��Ș_��	�sU�a�"�B�jF��o�Uq��I�S+m^�mv2	*�Z
��
����?�t�@���|Ƚ�:h��ڂ#{g���Su�^Z'��E�}��A)�E��Ny�k!�rh�x��8TT��4�	��cV*g�#���\�Z"E�L�-&�oq�z/6�w� C9�j��,�a��ƓR�w��&4�e/��sA��Q�lK��K���m�����TK��F:�#��{��]�Ǹ�J�!�tS����ڨ�v��Ć�mi�����g,�ߨ��k(�W3������k�цЬx�QZ:ʷ!㧂qoќs3r���A��,�6��)h衵�Ib�v�ٷI�F�P�C��&f\�1�6p)K}aF�a�����p�����.5�.�r�@'��ȋa�:����vl����(�3�U2T�]�d�1���0���`g;���@��ٍ3R�Z�Hk�����	��]�5`�'2��Kb�O�+��	���4' �V���o��yժVg�4-;��G�0�K�ަ���z�^yi1=�]�v@آ�^$i.�$*5e�b��S��I��)掵