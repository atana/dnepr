XlxV38EB    12a6     4a9�)�C�y¿vͷ��ȗNq?^�>]j}�k[����S���H����o�۠�� m/*h�0j�3��&n�4�c�/���o�vo�R	;R����f��"�"�A4�nE��"�z6�d�?`��G7���&I����+��K(�I�to�7	ꠠ7�`��3�(1Z���G��t��@3q�v�M䉧�n2��Q7�	���A�Z�()dn�e+�E�E���o��d"3�$הM�p3HH��v&�:z\��YM�<HץC0�)�٧Y���=���9�O�?��.�`c��?�P��h�=M�S�r�Y�%�͙xFQ�W y��C�=�p9�F���q�tT���W�����m�u�}u�P��o�V^*U����r��6�
����{DA|�/�Q�/�pn߷\����`��Iԃ���s�F���O�?��<4X����=�25�L�d똁Yy9��f	�`1�J��,���ч?%�|J1R��y�ͬ�c%і�2�1���� D�,��ӳ�"��&I����;���x��9iW���Xl&��IޱQ8Vɂ�[P[6�=g�"�p;&%1V�AW\sֈ����L^KB�Or&�\��3W���s����Z�($�W�z����@n���,��<�x�@b[o��&��J�t��8tj�Lh���g�n֟ǹ{vg����%F�����n�E�c��I����:�,E�@�L��T�:�����)�־�~�������u���a���p<ƻ�\ ��̩2 P��۠���o�({��i�Q��M�;��Y|hw2��9���L���v1��v�"&�M��{�@�:u�ߜ`k�m��&�ۉ'�{�ٕ;����.�]��gS��z��U2�AN��^�K.W}�� �ɗI���νlVD��/�5X\����z�X�W="��5B�6}m���dJף\'{0�R�h%!P<O�Q���7��\,���C�Rz^��y�g���i�4�h�k�w�w�`�@_�F�Ư��p(��;v_�aH�{�?�uY�nb0��K�ow6W�j;���u�莦+{�O���k�'�ܧp�0p苕�<PtVf��7h�p&;��ي�߄�JH�����{D~���]��#4:�x�9�a�̼�NS�l*˺�����)���V�lZ�"���!8l�:��cE�ŕ����