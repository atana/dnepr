XlxV38EB    202a     66d{�ӻI�U����3�3�Y�jDT퀂=�g�X�K,�;aʁ�z0֙V��&=$�,�,%�8�ّpi��#dJ�^D�o�-�\��sm�.�&l<\<�c2��:C��]:{�Q�0`���3��ŻD��R�!F�A�W֨f
T��:��y���C� K��_2���0��X�,��"ƕ(���=#aE�;�P�>@�*�vi��+ ��v�S��.YHڋ����m�Ǐ?,$��o���y��7F5j(�GГӛ��+����ۖ���Ҏu�k��(�4����=��1=K7G��Yb��
"�gf���$��0��ku�l�Yw:5�LO,�4�4*����%�&��d��W2�I�N�X�#n�]���7�9-\���������h��M�2�J��٧,k�	g��,�\�D�%8]v��=q{�W�a�Jwgb0�U�d~�����E��5�5�TRi��n�4�S~�Qy���x�uH{Ap������7����Va<�o�G�3�Ha�%�E^���5�qr.\�GCՋ����M�-����5���� x�[:N��[0!Љ���m�L�Z�/�e�1�+���6r�2�>��k�TŹ'JG�H��UY��j��W1g����9X16G{J����Bg�Ry^ݥ�H<�2e~�����2)a��2�|ԏ~�p�+�0��n�~X^� i^�4A�l1��X�4\�� ��Q�N�0�UC��LH���$��4���YY7�����A�\Ւ����}=_�rrx�r�5h<KA���Y@������m��A�T��"_����o�@��> @\Gg����*}C��9Iw��0�hoR�(�'�&Nf���F�F|*nAr���suC'�ݲcw�h;��'ERo:��O

��d����iݫ�F��y�xB��>�]3F6�Rt�F,�zZW��J[A�j���q����BR"���'B�����^p;��ϫ?�Tyk�A3�=7iU�U�?;�j���	�˝G����� z"Ӵ
���S��J��*�ἶ���M,�Ѻ"�jQ��i��_f�TA�_�%B=^ǡV3-:�G���w���n���^�=�q*F�|y�E3ٟZ}�0�84��"m#E�AN���75{^��g)؞r�$����m�@'K7�dSS�ɣGfq� �:~q'a���$��4D�wꗰQMxz�
^1?ŉ0�{�<�Qw�2���d�?OĮ[��ujYa�y���"����]���e���w%��D�B�uA���Q���$��y�M.�\��Yos��7�v��֨�]�L���v�i�q�V�aD�&h�����ׁ+������7W����A!�s��4�ST�Ŷ?�ld><��1���ԐvJdO+�Ő�*���Nd����DJ�;����B���*&�I�JS�Iia{_���keӾ���J�%�8kd_�h�t�hb��=$��k)���� ����q���>���-ѵH1|�����Z��9��q[��O=�J+��{]�6�������ד���M��	�46�D�i��Į%G�hLa�)x�[�F<�:h�I�S����������i��B-@	]�P�M@
���i��)�Xx���ha���93�u�˟�S�8C�b��xȜ.�