XlxV38EB    233d     8f2O'$�= XX�º�_0o�5LZ6�ȥd�/�K`�|�Q�J3ڣ�X����a� K��˚��.z�Y[{vL�G܀��Q���[H�zx����wZx��K*!C�O�����X��cȖ�%�{�C��ϟ�v���`y���Jg\sh4��҇�F
ߤ� ����}��I���E����x��e��S�KG�ؙ汖�پ�ߞ���i���=��!yP�?l�1�z�-�VԄJ�a�==��>�.b]�+�0�5P���W��gD���2�4��.1�ք�s��9o��DE��S[?r(�(�L�*�|���ԃ�#2_i�m��YS��7U�&��Q��!$��;���>���=�{t����9��L��l�\���9��UX��j����Ⱥ_ZR����k��j5`���ag�૎�93<��jh���79Nȫ;ڬ�G�����������U,��!��^�fY���ÅG�D.=�iᛇU~-��7އc[/BZ]�=n������9Xu�O� ���������m	�� <+�������Υ�G��>��Ƀ)/�=/��?���d������~������kCd`��$�H7�	$����Q�ª5Wd@���o*j�Yq|�����)����}:��hhaB-�L���z4�o��~�+��ɏT�v�����H8ꢦ�� ���<r=#�������L�3L� RS�����M? hY5�,ޕ��׃O/��i�r��s�l�c��e��Vv�"�����/Q�����¹��0�Q���VS\{�����-\�ª�~hQ�)��/��x���^�V�����XS�zoi14%t&�8p��Ր:41a����;�����A٥$�jb��t���5�l
zln�%�p  '�B���ʔ�b�e����m����(~�K�Z����Q�{0��bh+f���w�}�{Y���i���!i�{J#V�|=�,�z�v�f��
�4>0��������j��<g^ug�se4�f��i�M ��r��K}JA쏇}�f���l�yLE��x��&&7�-3��|��R�T����'���# 	��K8��j����ڼ^�������"J��m�O���4��V$r%s3ƺ(�%�񒣅O��8u��"��tU�
�[�\@k��������z]�]7�?S.�G��%#�Hz��G%�7[�v�5P���IQ�ܜ��C��o���Ǘ��R퓔+�,s��Ś���r>B���o�+FۦX��l�ӯ�':�!��.Z�y�d�N��bˉ/�Q�g�i��21���H����Gf�F3���I\24�N��9���Xl���hz7�X��Q�I5e�|���i�l�$[Yx��ɡQз�qbOƑ�D���{�FIKOr'��N�ћ�J�C>{���#�*8^11������E�������﹎?k��Lճ�����@q�CS�"�H�&G�N�����	.�E��dRO�h�;C�|Dc6e�98�n�ep�|4\�_`�X?��brL��.d��)�N2U�E�v�y��+�̊���`�/Z��6�o�G����0���4�4
j} ��S��9�[kT�{��r�n����;�U����F���0�+���FH�mE�XCUn^�a�!�Oh�(}�%�a�����m&p�l.�[c]�a�=wx��1��3w\r*p럢�*��|g��2`���ތ�B���)kE��Ȍ��Rg٘[�]��_~7�e�LWh��i2 �Q4���[s����2����C������b��T]�����	8]-��o++4����Nf����S)g{��,6�������� �G�B������ҪŦc�n���=4�\t�%BM!�=)�A�5 5�0e���1ٷ�R�L�ɓ�}��ږF�~�r)/9����M�{j�\��58�=���O�ʥ�<̊��̵�ë�VX�9%�X �s$XQ�̶~0s���!����e�ǧOw��L~BR�W=�A�I�ܱ:�jX�=ᕧ"7YȚ�?s�ĉM�baD0���l�`�zK|#qX��j3C;���͑�,�垫�gH��*.��\YA�Ɠ}(�Fx>�'m��So`�uس.B��a�<�9ڽ�5G$N~��ₗ�	ɔo�5���ُ�O��R���t�YK3K@<�X�km����IЩV���3B��w#��V1�x����2�B��Q��Λ��BmX��_=��9^�#0�Q�p���b��=�7
^