XlxV38EB    1c3f     641�8��!�� ��xW�*����b���*�����ǥ�6�'J�4%B�+l������7.�c�E�6��H��jP�4o��r�'Cq��ω�
�jk���le��(hT�(��L Wp��3з��
m�J�ڏ���[[e�6\�� �qNĦUĥ��2R�D'm�����0��t�	 d��s����:X9�,�*p�2Dx疈��q��w��l]��ܥ�E:����Q?~ ��W�(��W��Id�u|J8֌ԣ���1d�c�ؤ�w� R�ڀ�f������V�׆����J�y���Y�0tݵn�?����}�z����x+z���˪�ě3c��\<���$I�Z�յqEmVQ��A7�(�I���l�����\����wSs��H�z��"z�m��\{ŮZ���OA"`����#�cg�3���+�b�볪፫���7D Tb�2[.��2��E��Y�Փ ��(�;������<d��sd^y��aL��=Z�1f��w�"�*8����$S��v@��*�ſuu2���Ug�W�{�K�2���q�޽�1$�;�A-�V|�=[.uMtx����7��g��a�&��:��V�1��hăJ�^���y�%v�(~v
o�P��d9mON���� ��ۊۛG|]��`��DG�\ʰ�[�>nb��)�u���k�*LT#���|\���vF����Nڔ
 ��{A��3�N/ӏm���m�K{�����S�5=�iî/��D�[�>ۋ����̣!S�R�D��'q�:+d��?<�m�-����F����y��/b��)�K�(L����xu����C���������\�������^j����̞��*q�M�6�L\gz�'\XfG���� ��]���9яz{E�Amy;ӕ�6( D��)���'Adc�4�J��H�����|y�^uI�J@O(#�@���\ji��F%�P��SS�o'�l~�]a�  FG�t|tO�j�=�w�Z{�97���Z	j��ޛTx�i_,�ƿ�<P��LB���\�x�|D빻��S,��4���.v�[#{."�{���n�߮�d@��s��jt�A�]&Q�y�{a�7Q&���H��%D��J|��R������m�d�}�޺.��ؘl=���0����r�|�>�33����TE7����E(0S�Glh�`ݨp�4�K(�>(�B�B�rY�nae���xR�-A����=i���ɲw������,�F�;أ�ㄦف@�)�N�^`OB
w
�wfG���Uٮ̓��	蜛
�ڴο#�Re�m��+����}�f�WV��@|^w�D����4��I����j�+�+���'�"U��[{* d6���9C�`�E���tp���O��AN����)m��1o=z쪄s���(7|'r}�f�Yɑ&1����o��H��/�u��56��Jn��!`��f��&]��_�qn�� ��|/w�N��ȏ�'S�˻E2?��ݚ�i�d8͒�q��M4��wp˱��Y����2I�=����R>�2� �������<	��C&]���N_�u�w{Q\dW0#[Z