XlxV38EB    43a6     634~��E^�@�s�Y�$�!��ulh�A`TF�#l4�_�U�J���m��^&�X�׋� J�XI)`?6������	xV}Q����e�2q������`��܎�ύ�k�U���9 
P:��¨d������dk��#Q�|�T��Bt�*@���G�9�{�Gdo"e|�'����֘��Dāan���J'�սx���Q���X�'w��<��Dq��lzȂ�r*줆��(qĤ�}~����Ɲ ����Γ����B�*}��֘���k8/g=�O~��D�1ֻq�d����5��v�T!i>�#�No(Z2�А����Fq{���&Q3�a��b�r��OsO\k�I�W�&9�`_��Ey�JU3�� ��W�'T,�գ��]��v��꼗�٤�Ř⮽̀:{ �XcI��
�{��ռN�����5������>�}���xC����sZ^�}�Fw������)3(��T[�������y�D�S���hGDL�s�@a���j�~-Ά4�>�p��f�{x����̢Y��iIR��V&���� 4����<���m�#��}R�	�ł�����,K>��\=��H	6�P��~����,%̟��4ª[0
F׏�Gi�"r�qJ�5��C*�K�W7O����`1��cu	�->(0�9UlNL���?«F&Դ�&��Z�}�f�vOC��hr�]wD�����lK��T��^����b6\Q^�O��ce��]�wޅP}oorb��T.�H[���y�P�!���)���jĖٞ�Q��*��6�5/9��4kҺ?��a������r�#n�K>�D$nd�^�8='{<�VzN�w+�>��7v\
s긍�0�i�̀L����ZBz��F�D9X@ivvoM�� i�Yre�Qh�����.�� -�m��2+@��6�|��m��K=���S>]|����l�O�2�b>N�#$��U��k�MS�oa�u<�}�Ѥ9w��s�l��]����̮`����;85Vgh���:�]/��C��$Y����;�`����\.)��t����4�ʕ��Èb|�Җ�t��TWBl	r�\��FsjV���lgٲ��ß ��T% �kM��$5��[GXb+�p�4?d�=��e�������ʿ������J��_0f�0�����d<?�%�i��G@yO�p�w�LFSo��ScX���<%� -����s����J7;�FǤ�cB�m�Z��DX�Hr�)c��J;BcFU��ࡰY���y/x����'����?gr�q�ɾ Nv	E������+��2�#�'3a�t�^k�=��K�	�x}by��~uR*�r�$,N_���HT�a���;2��f�b��!��I@�W�Ī,�
+Duw��>�}`��,�X������@%+���z~˅�4�n�����ź��^�|�}p����}�~��N�&���:���^�̤��O�m�m�G�1JC�ڼ�� ��s���L��B1B޷���8N�G�UϷ�T�G,��f�!�����;�ٙ�ִI��)�U�`Sdo:��FW3�`;x��kd�	���+�