XlxV38EB    2ef8     a69p��{u��S��5��ypΰ��a%�A<�$�ږֱR���R��}�ddm�`��X�7�?~�s��/F{5�F�i�:��q3l��H��thVV����p�0yp�L��H�P&�G|q�<��%$����� �`�EGJ�A�i/��6�X�����*?��`u�l��R�B��V�4�`�����8��A�2o6��<�ϻ��W�����W�k���w����<���Z�tT�X_�3�ѩ��tTu��[�e�zH-�J���������cC۳���T}��
������Q9kh��\����2e�[�%�:��8<$��e������x@�b	ͅ2
�ׯs�-qjo���ٜYs|FD*^Ɓ�>6x�_%����t�N��s�m����R_#4ˇ9:�b�����4�X����_���Ng�$|��<��$Jόr�t)���ڝ���x������*��S��X«��bz��R�ē��������Q�Z��rn�(.x�QK��I&�����4�9��˩�j8��LW,���;�>���Q��Ŭ4gD�d�Cm4l '�)V�w�%��?�_%�G`T�'��[�,�l�f���h�e�1�{]�����~M]��Uu	�S��RU#�1�irt�ya�5���l�jq�~Q�q�z��?���U�D���PțllMQ�n��-�S�:��Us�kl����u3�ͪ�j��9sFWgǸ�50�O�u>8�3���튭�W,�D+h�ln{�M)5ڥ�<�5b���b�a�EB���-C�3���DW���pSW�uo�0Ii�����;<a����&��	�tRn>
��Ѧ���Y7�����]A���a���S/�����Ga����XeF���!0��=���rx���}WQV�1�����P=%7��E%z���d`x�����_���B�c�Ϲ�<)��p̾A�\�
���1x�*��,�+�U��P0o1.��������j�G�&˝f�U)��~��d��n�<n�(�@ׯ����a:��'}.m&tg��Ϥ݊,j���挌V�5�4�0���Ǡv����n������;�Z�!&��$���ӥ�'�s�"���V$�LW���t��!�ɤw�n��fžqh���K�r��ѳ�k+a_����:����6%��8qB_�	�o��^����^ԇW"IHY�ڄ��e�����4*���"Vp)`��D����d�$����W�2���j��+5R���U��:Ob}�rnCSr�-n��Ԯ�I�9 �(*Sw&��?<�����8����ɭ[�hv^k�u�5������a�z�E���	����jG����y�HW�l�~�2Z��b0���H�����d��b��4#�o�%C�/���7{�g&�A�SV�>��R�[z�#WM�nO��^F�](�x�����AZ�)-B+%����iEsޢ��娌�o�"&��f�z����LA<��bǞb�/�5R�mf ��U�ORh' ��L�Ǖ+��@��ʉ���m���D�R��`�'d�XR���ы�q3��uj(�N������m\^ðr�ĩ��;�h������Co�1Xː桸 �!A�J`�\����Lٯ�@�-[�oh	�Cr�7��^��zS�#��8���T������%��Ħ)+���7[q�68n�3�[�0<���$��~��bb"�If
����S)߭x4/%�+|�A_B�A��`��·�p�P�:�HŜ�f�1.��Za�aI�:�O��i��K�}��ǳ�V�gmҿ"������3!�M"�t��������DKφ/G�Od����lD�O.3UC��Y�^[�}�׮M�H�w;
�6K
���w�Ћ��A��b9(�W��@T*�����	yY̕ʎ�]�Fa5"���ho���4D&��,j*�i�o���K|�#����}߅A��d�e�%G3�}9�['7_��ѻƂt�n��cU�'\�AS�
��hZM�=#������/M�2M����8Cbi���>��b�z���6� �$Av�~�;���2^tOZ�~�9�����Ƨ��v=I���h����Ӟ�
0P�x��%��P@=�ϴ+�P�}F��|��Kϲf�Yz�5���񓥏3���(v""�$��H�8�ֲ���*a���|#�bI�D��ʓz���w�p[�A_�+�o�r� ��u���"Z+�Z��:�mm���O�{MW%0��qɴ�)V$���)ŉ�{�M*�c4�еe�׎u	_��SS˫5��Ҝ���P2��)VRb�'�G}�W���@��%��'|��}��V�k�m���qV��\q�����*ܲ|d�w����XpCJ#?�߃���P`.i�#��п�i��R�����)�Q�>���v��r%6Q�b&�\���J�=����A����ͱe5�%��w#鸽��"�%)��<��������:s�Yո��#�"rn_�l�l��@�q�=�1P��IĢ��YY�o� �tLԛ���F{�B_��{���2�5��/&%�v�S׎���������n~���{��8�x�Y�ND�W�|��}�����R��oJ�I�K����.
��~�(�ϔ�