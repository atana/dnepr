XlxV38EB    1393     505���
�)�I��=��o�Z�K���-���+T>ؙ�ڗ<�E���2�
 RM�B�����4��6�跛<���������}q��Yt\��*��B���5��ތ^Q^�2��P+5�{��lU�Kڹƿ3��y�5%yQN�[�G�u@g�zmØ���Wt����r^îM%����*庼��nӯ��RC�9Q5+ՠ�����7��Nb��R�Я��8CȌ�i����Q�Q��V�K�$�Z��(��<޶�&g	��)̗±v�y��7P��t��.<�_m���r�����o�������?:�b������̂�g̯ `�L9H��x=d�K4���91��=�����ξ� �2���f�]��"��i�|L��܍�*�l��߅!�Ȫx���mBH/Tj�S��A��`:%_�
�=Z���9��w�A!��~ڮ�=6�	���g��lU�����9x$X:�X����1ۃ�*�OS�'Q8���Tlz�T��
��5T�:~�~$f���K�)>3�f�-Oq�;�Ɓ]pѣ|*9)p�h���ʸmkt����.G� �`��phQ���H�B����xC�Φ�g>֡eEAT�����m�Ni�� �8.tU��Ҫ�_ fe����-��ZI����٪(C�$���2��=!�!�Y�6ڏ7 et��� f�Z4;��4��W�U����[�O�8�ـI(��s�K��*fZ�W�L�pk5�_T:w�Vg�W��$V����靸R�Mq�R5*�@?ْ(,�:~����� ���S�� �~�h\U���6�H��׋T P� �Pv���T	��f��	�p����#k!�f���l���׼T��݋
4�JH:�K�gl@zK�pZ�/��YR�p$�Yiߴ[��Nc��� ��6xQ����F��0�މ�N�����<��݊-�pH�[H����n���}t��fkg�!�`�����Dz����&&�ǐ˥կy���h����9��d���a	�0�+j糂ƿ���?C:C�"�'ue�'#���^��G���<�aFf��Q Ɔ`r�p���p8ى�}� �W���:��Bfͤ�9��p/ｦ� ��يE����s�Y /�ت�����'����r`��U6�h�h2Dt�m+�·L�ӑ�H��Я׻�]GB#%�F�|��y[�EL=��;�(0\E���#*�;�u�q��Ѻl� � ���Nh���u��#�`�����:����