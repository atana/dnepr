XlxV38EB    edfa    2118ϐ8�3���H�� ��~axˈ�l��Y�U:�a=���ҸB��ۜ��`����^�u0_?�E7zF �atX�>��WڜLY[������I���ֱU���0C~|j>����8Ph\�K��&�
�m��z"k~�6עޮ���7殅<)Ö&D[E�������>԰ZD�F�:�����<p��=�`2�9#sa~f�y�$�b���SZ������5B��A���LV�.!�r0b/8n��a��!��hc�x�ìg��i.S�[7ŏ���ͬ��(e7b�.�,�#�Jjf� �tj3^��($��D����z�A-����N��4�m��*�1��z���L,Eʳ\�'K����k�1{/��v�n�����6��F[�[X��Ik%w�OD�M��s~����t����M����"3_No~��ߗ��A�R	�`�Ҟe�P�?��oB�cv��w����aw���48D;�#�l��T���������\v�rGN�Fw�X�!�s-B�4��/ �[RB��PK^P���m�|S���`Uâ�mS6�m)�3��T�խ�d�#�p#��#<�e��|�>7U2�qv=��;?��1k��W����?�P[��0�}�t� �V����Q�Fp���yF��K��֓�e�?ia؟�j�E]��^p�<��+�w�6s3�JX����{�^!�.d���hov>��R��0��A�CZ^
�����NS������H�'�e���$�I	��k�]��_<���3ra�'
 ��9�_K�V����H	�h��}��N�'�?����x�ٿC�IE�3΂}���7�qRR>�ʣ�¦5D�O�um�c�%^���ď��u��>���~{����rW4��p��w�Dh��wn�b�_o�U��'�s������e�=��Y�����+�s�_���iQ�d<:��i�H��._�piv��!�:'�S��uw6	6"���ۜ���pϧn�p��Mg�ƪх��A.��DN�{��(k��O$G@PBsY���:�(�%����-�k�� gjkxH;#?���{W�f�Lr��5��ֈ��W�%���B�ֱE4*�B`o��=�Q>�/$t�E"2��������?�HF�1�-}u'�?4�h�K4js��.CFbi1��Ӈ��d�O���ǃ��}WSy���ܓbY�<��muv*ҙeT�'Tt�ADV;�U(�m����:��%�K��Y�O4���P�m�̫|/+��6K��
'���7^�V�g�x֯��-)�7G�p{!^g�.�Ε*�#�%�-q�����������֊E��֊ OqG�̍"�u�jւ�Jט5T�Q�uI�"����^��4�Fq�qW�wC�3��F�^�2p#��L�ɨq�����R�k"��`�c/(��*,
����0I #��9Q����s�߲�/���IIe�u	OCUhKE,&h:�!<��'�Gv߻��PC�r���˹aM�!�'��ͨ:O�k�U�v��FJw]0|�2��ף�����v�������.r�u۰ɻ�Dچ@Z���x�l���%yF���^ǃ�20�kP�d����3����#䄄����P�&�y�W��T���I���%H�ĺ�v_^-���_M�������S�(w�<�PN}�Y/����r��:�.8V��<fcg�*v�����$d9���$�a���`�~֫n���+ܰe������\�M4:z��N(r���ɞ�&�FR�֒S�z�uaD�V�9X�	yi�yo���D_��>r=u��q��@
��?b��w�rm����c��9W�%��=4-�u�#���4z�[���M��N�QG�}4{��!��^5�,�.4�!���@F#�����|�f�2�����XJ��e�$�W=a�B�v�	�!Iz�<f������ۉ+�*Aj��l�|�?0����$Tв��^u%4��ပ��>�0��B]-?�����(��PId����eH��;�����横Q�#]u�8y��R%D�bd?l%>JdS��M����1�{�:-�	��F��s�Uuǵ���A�����s����[i���L{y��C��9˓�H��Ú=���e��= ��a�oliq/"�2T�.A�\�a��u+}e�b��+,�чh"Q1U�ĀA���G�����:;�|��5�NԞ;��np|�$���H�y'h�Ĵ�/�b��H2���eO��"����-آ�ؓ~?�H��z^+h��t�Ͻ��Z��S{Y�XYX��1t�����!�!�þ�D)����K}��k�s��2����H^����s_�&�ΐSe�"�U��A��,�����Xxcw��غ<� ��w�6�9sՎ�ur;w;k�آ��'�IN�t�2�j�[x�[����,�@��~��('i}H���_���yI�&���-���C��|sS7���urc�N�PT��&���������	\(sN���d�;w{L���;��}=$�dIV��T(�Ȉ{;=�w���{Y��+�o[=x���E������4/��]b�å4���Lq��]c�Vp�o����r���s6&t,�]�M7d�.�4�(�?]:�WG�!�s�J�ʺ�Z�6|�aAjЎE��)�q�V3�d��F���ͨ�B�`���O~RNN0=T� !ؒ���17��^�H���Ŗ?s-�D=}xy�Q�(~^��5�nj_"��3/�Ż�`����H��tS�p�Gj�R�Jffw�'��~ܥH���I8�V�n�8���}Փ�{E�fOC�KP��d�.���ρ�!a�U���L�_	8U����:D�,y�)�3R%v���^)���)_w�ׂ>�/b�5�Q�4}�5�oFsvz�Z��vP�2�c1g�0m3=��(�a�����?�L���N��&c�w�nN�Z�c���^m�B1l��c���B�Ľ�3ʛ�z�>K]�;���xU�O��J4�a�6��?�z,a_7���	W��ʄ�T#(21�^�8�H�����%�b��b�/+E!���d{���/�@r��Ai��5�ڃ������~Ivzhra��6�!���P;i��<�+��$���k��[��G�K����B>�W�OӀ-�E����:�X��՜S�A]_�-D]@�dۘ��hH�@/��ò����5R��{��Q�.O�D�V��[*q��H�;َ�]�r�F�c	b�Þ�g�G�(��e��n�(}!O
�Q������5�L�DXЦܴ�U�"��ʁ���w�Y:�E��o��_���β�t:���J��x]�?���5���ۡ�K(Σ��^��ݷ=��["X8)��wn���� abu�������o-.I�דDvJS
�8�����J`]n�pG���Rם s�b��*b��t4�Z%���i�vD�~"�����Bj::��P����u���@X1G�P� U#��Ä�5��r�T�9_��D0l��$9ʏ���q	 ��:4�⊄�u@Ǟ����iqRcX/1F�mM-UӦS��D)��2 NN�=*#����W[|M����h�ԏqV���(���sK�/S��C�N�j�@�֢���U�-����/3e�>�O�/Ԯ�}s�t"���L�JOc������OV���7�k�3*�,�~d�:Y3�ӛ��O;T8�[����p����mԼ-����,�n��h}1�	��ˀh�MX�v�扐��ۇ%�)gB��w�%(�
�Q��x�R�C��6� ��ԞQ��Q{f|m6�(cs.1(��AJ=ه<b���ֵ���S�%�&UDg�JD�96��Wf�>�.������W���B-��uI����fOW�7�ܗ�A�h\��}�M
hߚ~���ۢO���j�ˌ�QI��#8s�CE�Q�ϼ�	��ò��;bxrG����oLͬ�k���Ug
��O�;1ӣ3ҵXY���iY�r�+�w~����~n/�ۜ�l���h�D>���W��Nµ&,̹/��+�gmu�z�P	42�i,�x��9��Mr�i�G��7�2/�JN��"[}ò�W�ΫS�N��FB�dH϶C�n�
$�$��T�c�ֳ���6G�A?���W%��#��V�#��s[�/5DiE@%X�"B82���Fd�B�Q��B���d>�13"T��ż�A��%8��8����L���FM�NV��*	>w�'�:�L2�F�xu榜�ŗ(Wu%v=1X��ŀQ^J�I�o�fN�,d�i���9��Y΍a�ɣ,��6v�_RMل>���m��U|{9�W�̽PQ.�2�ޝ�р�j����8�Ke�����)���1;0y8j�Q����]�.��o����f��4��$I|��j�0W��ԕL�Q�;y�L11V�m�D:V��7cM��O�߉@�qo���y��;ٶ��S��D�+r��@��d�:�?cP����O")~5�&h��!a�m�\���U(1����5��su8	6�������i�(0uJ�htG}��&�Na��;b5ȡ>ո���hy�_̲Ԃ#[��Pk�u��;��2�D�0ҘO\;u�#�}�b�3^�GQw��g$�s'�O������SŠ�ߧ!���!�#�r�}�X�,�_K´���#ѩ��.W��(��j�-�����I���3� �]�C1��G�!�݃�/�)*l�߁�%�����j=�ĨG&c<���Y�_!@�O�3���O~K:��i�"�)�
�;���}."�^�������a�x�r����A!9��x�3�������ޥ�0r��hk�1|�ڔ�Y�i����;�sʽ������ʀv,XEB��г�����ky_��Eߞ����&y�miX� ��_[:M�
�6�l �{*;�d8��x�aK�rn�J޳�U�F�*�{�8RˬeͣtFF��sc���d�g�xn;��e��I�9�F���ǁ�[^��aEL��ѭ|�=���N>�ױA�z���^XB�sd�Z���EE��)Ɏ{�qS�)�t�u���m],���U��=�dLa�_+����-\��';�5��5�/̂Cr�<N ���f�6�X��y�$��4ݳݢ[]E��u$e6����Ǹ��$;��J=D3	XM�q/s��Ȩd@�󒾼�d=��>���oV2g��iP���S�t����
7F�be!�9B��|Hh�����t�� o�2�[ƛ��0tWl������q�JNi��)&{���q�9u6:d��0����(���7cւ�13oNv-��GQ�m�9S!��<�XR���TT�|���]++�|��Q�'��q�@O�:$j�_�e��挶�(�듪b�� Ȩ���òWA�����b ��V����̤�hfk|�:�|�|D-����/+%�9\�^*F~p��#��է[d�u�On#2jE���:���Ȕ��f�dP��c,Ǘ���)JǸcE/6�.{W���#���2&C��GY:�_\Q�ﳣ$�IZj�+�|��e;8�^;�=	-7G�ӋCj)*�3����K&�DY�����C�	f��C��@⻹<�q�x�������q�����Վ��H�kF���[�ǥ��B(��&�.M�͢�b REp�ꄉo�X������B}h�c�OӲ���NY�J�g��ӫ��	(����О�� J��՝���91���_~p�L!���ݺ��Gu��v�0���v@��$�h�6P��[4��+Z���5S�-�<\7ڟ��C}e�Y}#����L�lF�7w��=_0� А�����\��ޤ�Bl�W�k18������H� �����E��ߋo`��2�{D����N��V�@��u)�(}$r�(s��@��2�G��E��(Y��Я���UE�����@�����BaB�~��
�M�*b�
���G&y�&>_B�]��& �RY6W�F�e�T�7���\��%�O'���e���%��`����L/���%�aCu�������|6�DtS$���D�[�����>��~y).ϛ¬ e��U�t���Hj:��䥘Bi�#�
�}�S3oxֈ�� ��dT$�/���W� ���|:?�w|n��'��W�p���yDK��� ܷ_��Q���b�ht��?�Q�sʩ�A��:R^�R1r3і��e^�ZzG�8�	���!ɿ%�/ �1�ӏ�{~�xU�f��i~��$��)���s�Q픒�A7����:���[B���X�Q�O��(>`�dI2dS��|H��nϪ���lB����؈:U�E�I�lT��b�_-��:L�r�I���a|�t*I�ƌBu����79 ;��o�*�Q�) �G��1sm�d�=��l�������p��R#pN��ި�����{��W^U?T��D�1�D��h�Eڤ@�5p��6�$����`�zHD�xڪ�C�$b?����>�\)��I[<`�:E� Jd��>����]z^��-�Z�^�]��ظl�{/qaN�A�+I�5���xa��.�8�/�:Β���s��ΦW��w�MS��~fu��~���uy�됰Gn��*�W�b��^��WT��$'p�b|*�Z�l���+.>i��ص��18E�j�s����C�j���4�!�T�&�����Ei<���ta�TG4Y<>Y�H�!�&M޷�؋��2��2M"�����x��U�5����ƃ:�<ھ!���+��oa��V5����Jm��{�C��C1e��@m�{�I��3�#�"��jR��|�	ΌG��	xp��@�M�(o6�;�F��m�[a�+�f���܊�u��(��}0B�c���udN�f�r-�j�T_�Z�ly����c�wu�Z���˩�*�e"'	�yĤ�����:�G��[�o]k���S<(5V��nU��w�����9������Ҧ�Eʓ�s���o�t�hԓz�vn�W:�q����ڨ�.�M�X��W���Y0�	=�w���GX��ZNz��y�s�������,jrb�9�&̃�qin�}�d�S��V�nEk�$������H JWk�gKҼ��/�wZ�ׅ_�9�=��5 ��a��<��S���=/���m,A�;>��{�U7���y���g
C��Ĉm$���I\^�A����G�SR�1pQ5����̎��Z��5�Bdr��(�(���|�C�~<_��,���V�\ x�	��i3�kip�#jp�������_��%霌[I����-.�J>VsP�qQe؎u���LL8A��a.b|T����cZ�K��n�>������#L�K�\[jպ��](�"���k� t��v1q5��!<��l�!��}��$�$�5LaWv�#�@Z&Wi��!A�����[���(��}Ĵ��~��ۮ��r!���W.Ef�����;S+jY�p��P�[��P�e�Xő���e��'����>!s�c����WP�d���kX1!��*��({����ߚ�\n\����8����ED��b��|�MP�_Q-�J������}h�G%G�(R6�Xcu�����(`-�r�v���Jp��x�x3wF�meK4�3J�K7�I~��K
��)���� ���P ��v�i�<�ˏ�~�K����=J�T����4;F�����<	���kj8�+7D��3zԇ��?�Q!˰ݛCx�(/"�[���l�a҅;К����LaLڽ�8v��6���Mz��Y��~��7\���|k^��&�:2��b�)��rc�{��W�T�K��7�!���r[��\��I�����~�q��@���4����1.nQm�PB�|�ɏ���5i�7����F���LLBR>	G��/&���`#6�m�-�jY������g��.U��@>W�N����)�O�������,���X*����ML�9� 3�h6�W��y��a�X���lY�.q�!�#h���\�-���G�? �.W��r��+*�:n��f&i�%�t��z�f�e���Fcs��?���,��q	��ݎX�VR�
��8I�x1���
ľ0fP��X�j�S���%��B��=�	�dB)t�W�+V	�B��D�a���R�I�=�x�s��2��#{��sW,�y� ��}���W�G��oU�*��;
�G �%c�T��%ՕCMI�t�� �ȼlS}V�C(V3�{��%8����m�è��8�k��`�}����PN����%#gT��9!��!X���S�W�����H�]��`Uj�