XlxV38EB    9b1b    1978{d���O|$\�T1�$��.Wt�@�\d���Q�5)��
`2N+���6Wơ[Q܉�1��K�rs�����^��z$��چר��NgP�J���׸b�E䒡�|�9��N�����"��뉖�u���t�v����9���l_��z�H�l������y�
ti�^��&���F�_5MWP�e�4�˗舞F�a�cF�k�I�hP��s�,���%��-�˫E��>.���$�Oo�#�{��Q��hPFR�$�[�>��<*�9�^@ӜNO���p�=�fHl����GBL�B�ꄢ:��OėO�H���Nź���n�a��4��� E��
��n�s�bs:B�M�aeX����|6
�s�ۑ�*]|a���� �k�/�k�8���J�˟}b	"di3��yBȊ)ڸ�:�ZX� ��fec[p����v�7���7�5z�8��Z����m.�+��D������ܨ��������ˀ�g�`�A���&>�����Dv�V�J��C��r�ڗ�BnV�����f
��ZԢ�;B��}-e�a�o'W�ςw|�U�6ҎD�ʠ�!-S�s.k)3�>64ǰ�.M�$ө4�$(�,�j��0�֘�Uu�KU�5u����U���ɘ��@��Ѩ*u'4�M/"l�� ʴ �]�AU+˃ұO��5�yoo���<��q�(o��B���]=�òM3_%o�$G`6��� ��uI�0,$�L�BAJ�6p;���`u�7
��~Dؚ=���@�x�
����觐6�x
`����Q1S���$����O,��*�~'}JZ�Uʓ����h���+��w	81ɝ��M�m��\�0�H	8�Ի��`������6�
3���У�9(���k��)eG����a�]�JE�6��n.��
8w��ʹ~BD�6Su�Oo`aMm��]%FG�n��W{^ U3-�I�T�pS��B��ծ]\6��Y�k���e�%2��,��\p�1OBӄ����4�+��]��=���KO�b� R�}~�zD�{<m��|�+(�_GB��1)XB��	Z�53[Z����c�g�W���U֝ʴĒ`����3�=ٿ	E��D�w3��^ɏ�Z5d��v�h%�	�5@�Э�M9&���Ey�wZζ�ז��$!��̖�Q<Wm%WL���S3�Θ�#V�'9��"ȝSOf�Jw��*��5�����J��(�j5�;n(�Yd�����IGh�a ���aPW�Z�%M��_�'S
���e��`�|& �)�rg��}�������$Z�+A8Py(��A����r�u�*�c�S���s���y�K$�Ń�IfZ�%xs��Ơ�0b~�'�x�>ccmTȫ�k�|���B��n�r��h�r�\������p�Z2�t�^h'Cuw���(>���s�
����2�<Am~���f3�VQ��o�5�|���"S������14{D���ݿ�ԃ70��I�s�c��΢T7M��Q�i��SV�ۊ�%�z񲔯�mN�aoJx<$Z����(��X.X���H^w����5$e��ܤ�bz'�(�#��m@�2��TN&���(۫��ET��ب��];C�k�Su� �2���K�Uz�>doC���
�Dw���}��L��xϕ�k����6G��Rd4,��hh�Wu`��;�զBm�ˏU���1F��BA���-����k�`��{��K\v�?Cu}��S0A�I�_PP~0�Bɹ�|�iQT���_����6`�o���f����y����ci���չJ�fĕm���g�8yw߰Զ8�B�� S�J>��j�������c��f��[M�4lc�6��;'�#!H��������/ڱ�������p�50�;6���eq��w�{8(����jr�����Yy09�e;ŗ!pm�~|A��=f\����F�V'����e�F�����9J~3��pH����j���dt,W]��k�{;�򄢤׼��t���%�\�;�=��Vۼqi`$�i(�F���o�~������plm��bj�fH��N]+���z�q<��W�w#(g�xe�#�>+y�v�p�]��%������:T��n��ƈ��<��=��d�g�N\zF�ǃI�-����0Y�9���U�Dg�MeM
Bʸp�A��n�H4bkk&1K��yCˇ���@;���߈�mb&$�I��r%x'ZiY�}Ax��SW�V!���1�!��؇�o��Ů[?s ��dR���� �yPe�J��#�%Pn��ѧRN�6�E޺��K�A�:tx��X�^/��*�)��h^���\w��D}B����E��B�)N��pW��+��k������lÒA��v$>_/
�u����LEs��$�2���7�hv�a�v}M1ļF�%ϗU���v�:��f�="��d�w�HA�5���VK;�x[l�Ӭ�^�i���4V�è|�8�aD'�yt^�ɂ�/�Ռ�c���d�v�����bh+?CrT�nU��{f��ɧG�eof4K�{˄]������k��"��o�}Y�x�ĚZn��V��L��V��͹�~̜6#�*�K(X��Y��;{GՔb���e��E�d~{�d엓�T_���Ht	����RL�x��[z���*KLhT�ulɦ�o���$0��%M�%��2.0��u����n�ْ�j-:?|�_�+oU��O�{�ۀF���	��{׊<Ѣ0(���Dh%��-�=+��r�����$�E�*�Fr����l��F_"vH|�_D��OԔf�_���y|���0���q���b�T}(���7]�6~�*����'Ŋ�܄�o7��a��/Z.�Y�/������r�P�0 ���:k��ܡ�A�V1����'��Qkl��=G����FfX~l-�]��\J3�w6S�@6�:�oQLé�����Q�h�x�c�p�h����hP�����_j�%�$K3$�`e9�H�`��}}3�!�B���6S�$�s��������?�,`�#�d��c����Q�)L��U�v$��鼃���M{����~��kP�7h�U�9b��$r�u�Z�A�"�^o�4�*�Gͳqo�Jx��H�=��z��$�q��\�@h��/}��n�|���	�Y3h����9���c�g��Xݹݒa���ZvD��+J"�rV�Y��AI:I3��>mM�EÕ�6�T��#��U���� �[n���(�-1�jgk�����06#�s;ٷ����4od�f��2�l�+I>z��Z��w�iH؅�r�dvo$��0��7��>=��s��������K4={:��R+DZ�N�(��\iSf�Z7h��BXoH�X7�TB�aN�����X3I��Zr�ԙ�L�!Yx��>$ܠy�r��ψ@D����9/�SD��-<��%��k9����i��Ja:��Lln�RԾj��m���-[����RkRu7ܑ[u6I�Z�i�N7�7�cB�ה��"8򴯿���H��b�����5�˺˺Q�P�}�<��V4
���l
C ��HT������8���>$.u��׼�)U��P$cF+_$���R=��� 3�f~�k8ɐ���"���8Ȧ�3ʠ�N'�O���%G�[�q��:�d��Oˢ�t|�?��On}��HKDh� �W.I53����,<EHA�P�V�I�E-�VFR�g�C��Y|��,�����H�ϯ���Z�dt�����
��\�gZ��3���������9��x���.�rs�a�q]+�Mz�8�,��-qZ�Z�
�^T�^P��q��?�|��c�3�S�!1J�%���Z�@�^��Ztl�
��4)f;P�P�������l��>�ތ��E�΋j�ÆE}��q�ĺ�11��g#��u-b�́�/|ڥ�.ȡ�a
�=^��K��NP^�ī�R��D�����/���^�U#�n4٬.`0!��������v�
xr��+;(\�ȫ+�\�����m�u���g��#����P�.6=��C��FP���a�2�Dl�1�P�uj���]���JB�j+=n�/��][��73�W����t\U�܉R�~�����a��6�j�/;^��'3"��]s{$	��� ��ʫF o����[d,M�l'����d�� �D�Xq'Ux���4�]> �O?�W1�e��:����Y�{�� sP#�9�r�Llc>��4���eƓDkpb�	M�����l�3�6�KX�\��G��LMej?5��h���.Ҩʏ@���g� ���t��x�p>����Zp�YOo-�ڪ�5�uC0 ��� =NݐX#h����Y��$4��1�{�J����;��sc��k\g(�[OPb��r-�^g@��:m��ҿ+��_r��u�i�#]6Fn
,D��?��G��d�M��N���^�qZ!�0깴r���W8i¢$G\�]Lc��l썢��Wݰ;�S>��>\�܈�gdBJ�_��>�{�Ϲ���n��S@��$�4��lU�thX����m'��8pv.>�)���mrO��Y���g�l�8�����tt^��I�$�:P����a�4y@� �@$śW,^��ɘ�{N�Q�<^�y��`�)���h��+NVJ�V��������Q�㞭ory��nuD��K��/ւ��W�3%3�'�2uA&�X|�QE�������.L?���k'�n��~��ֲx�0�MbH���.o�M��/�x��]��ь(g0H���N��ul���&BB���l�����B
�����ϐ 0x99���vÅ��a���9�j�u%�%�)w����e��*�'���A�;�#���|썏���u=(�S/z��</���84_��o��^Q��`���`3�,
�g��?��K~�$�~h�?X��&hD��l���U�X���'��6���'��Ej�>����p�������jA,�{" �-,O��L�R��A���̤�ۦ�d�7�����m���l\4U_���Y�0�_+]�1�����p7h����f���{�A^��@O�"���q�*����t���bbe�{GZ~���6js95}�������L�Z>X�����.���΀��S�P%�#:�,�J�=PJ��&��V� 6�y��f�V_#E�ђ	(�:Z�+�O�%��CC�1ΦJ%̿y�8�=^�����[Ew.1 ]��_�e��haAL]<�W�ʞ������U�K2VBZ4�����Y��?;?`6�&�ia�BZ���U���޴�����*�w�N�_�O�~Y����ˏˑ���Ȋ*��9S�N�^x��@QK&J@��<�,z�`e�U����3���݅�;���S�|�J����
^���<
�rk�LTn�6��=���8�E�m����k��)Tsxo��H���\|�H�\zN�O����9k3�X����7gDh�^����??�%��n�+M����<br^W���K~�����G,�ӌP��46�a�nsߔd���{�6���3pN�(��*_B�y�U�9٤:Q�����0�a|�K��@�H
p�-���\�����:"&c�"�^�9T}�?���M1��G��QMw����)NrɈ����@R�����C��ȂkF�=�]],O0�b\R&a}�n�DL�M(�A��8}D�J�~,�S�}���^�=}��,VC�z�'J)�n�C.H3�XG�..�b�Z;܏�M
�{Rz?�:gK(�_��*h�La��'��qSJ2��{�	L�u?ԴzV�7Ѝ�>O�l���f���-LQ9�C��<,8[�Q�t�2K�u� Z�Q��[��&<�?0�t:|�hR}��v�=`�Ϛ��L����G�:�4��b��`r�,����g�7���W�E��~��
�{g�`�>�=#�q�.XF����Xd��gx?Oddח�p��ۆ*���o��X���� oHQ�:nW2�*ѳH�#6W��g���/������g���+}�%�(��@��D�#SX�o�;y	&�l�0*��o�7~���P�^Lf^m
�5�U�M�8����'���WR_c�b^y�����s%�1�z��#� �c÷�!�2l���R�ko��7���N��=NE3�<f�3_��~��S�ۯG%Rȇm �5i0�x�p����	��Vz�Ր�������Q�ץ	�0�>e��P[N�%�� ��@��z}�� #�åW���<'#z���
���A��n3x�q3�i�s��ڬ����z�����P���͟�O�/�u�*樳�hr��j��z�׳��^� <X��t��+���z2�'�$9(W��|P��a�f��-��	���G�/�@�Y�d3�F.��X�ԥ���j�}"���qݘ�0�/��Sv������ӟKj�?�E{0��Ye���,�����8�#,��;��