XlxV38EB    1302     52e�W�Y�-��}�(@��ī�_r��3�|W��vau�z��A}��.��
��̎�
���bx��.�!�gd=.*Q����0u�cF.��{]�=@�o�*��ZkFKyW�g�Ak  Ta�zĤj��i����>�����i�8�@����3�%FRh����V��jF#�.H�N��ٸ�Ko�ځ#U�6��<^���5��$���w�~Y�g�
�𽄛��*���e���^��6�G3�-w�?5��t��>�f�_|�o�����ASC��Q�r�D�>������'�;K*vji�[s���Hn4�n۞���Wh/�c0���-E�Q�?�
�*�OV��|�8����I�]��S�K��N������uhΣ�u0IU]>c�p*ųvJ-;�D�Hp�.���s���[��7[	4)@ձ�>�kt�%P�a�1��6�\����σb������S�b�� *��I���*�싅��O� y
9���=�,l1|�u#�/$Ħ������]�Љ�����J��ߧ��O��W]�8"���+D�yZ�����O�o��9��#�n!Hl	@�3��݇y��Q�Ԙ�}gO^�әg���Wʸk�J�]uZ+8*K����������_=���V�uBi7�8���3<�
���b9�O���=�hC�
*�2Bs�'k>Y��ƁP�@��k��Q�J㝡d�F����	]8#J���o���1ނw�ef�)qؾ��Gv���aۃ�TK(��vW�uʮ�_/�"&�P��' ے:u1�*�riF!�Ma�0v����4���"phO���Cj��v�tk�Z�`0��z) ��P���궾�0]�԰ɨ�5kj�&|_|q̧�X0�B��"D<ڱ��8N��R��p�+BAJ�}�fq�3S�ۗ�c�iAF��3h"�C�t4%SA�Y��^�����q��0 Y���<?h��^��;kQ���0�X��M��%=��;�$ͳb��ks8Hi�3L����BT�P6P��7o�<Ǡ�@���+����{"�����c��?cq�u��|�͐ܵ��ԝn_C������fb�}����������sk��6��"̿�j�3T!Ĕ:� &��9�l]ζk����u�fgε��?4|���wrn�m�\���ÒVh"Yd���$��|�{����K�hw���F���Uu#h�I��`�<�����(L�G�~������V�h9�j�+�u߷kn����%��^hu�Ѿ�)|;q�
�1��U��\�d���Ϧ��De��?K���