XlxV38EB    327f     961�ēdEY�7$�n�D�tw#W�aX�)� �wY>in�Km�''Ʌ+�����E��੏�	�%�0�Rj�&%�v#B�^D�x�
�b����`�Hp�1(6�y2������b���V���M'fd��	D�����Y�jПz]��+q�zG<ͭ�AP��;�=Sx*��o2�D;�Q�p2o^�
�?���óB����y�K4J\Nb��|����Q�9}��d�5Ur)�^�z�g�MGJ~�=�J�(����T+�4ڽz���r�]�l������{�+i�x������� iG�Ǜ߬ݵe�tM]����2��n�_�um^]A�[��h'��W��?���w^G��m����vN:Z/*�$�"����b�$sՠ������@�K����I��y����d����*��VJ�j�քtБ ���C�s��6��Vsd��]��W03���M��ۗK|�Zd[|BY��}��������p�/�w���=�a�f�	��%�<�h�YB����Fr��U2�ܟb|�¯�ڋ!):$��c���z�(����Q�G�Ws�HWzֺ}D�%?v'�O�|���
���0O��&�)�S�3s<$��:�P����)���������l�5����U�S��)������U����@�O���[
h�����/VK�r���OƽX�i"�q�az�?>�
u{S4{�����԰�+mXN���+J��������cqojF��Ժ�@��x���U���T�H/��eCui�V|���W�����t�4<�b���	j��*�L��v�A��)�-��IG����miPEq�5ӏ�,?��W��}���p61�^ORTS��Q�)x&O'��! g�B�4~0���+�$�l,d#ҿ��0�.4���y78���nV�'G�{�Ak+koڼJL-���������|�����-���֤��L���sw���Y�|x��G��y���^��fhv�TQ�tkP�*�F4�nɽ4�2����ڔ��UC�|q���`�Lz�C�`�� �h�-�;mcX,�G��g�F�C�|.%�"��2�m~��[�I�m�
"\D�_�����?��v�J@"�䴰���Z�	���9/0~I�2���sd����d�@��焝
{� ����,{.=��x��|P��,����
_�Ԗ܁�P�}�Ҷk}��Ř
5���Μ:����A�jvF?�O��YL���Gk� o��V�� ���γ�o��-6Z�Yk�\����Ԥ��}`/�&�[���{B���@곉�J����qcȬ��>ۄL0�ڿ4��F:Ѩ![��.�9@MΤ%��0�������7�Z��+�50mK�9�$�,�a{��a���A[)�4�m�'a��XDTUG���
�����y��Lp��*�^4}�`$�sʪ��͑q������ߩ����N�S��#����%`���[��+����~>,�k���!��ϕ��^���F���}�S><�n�搣�`d.�c��X��}H�mX�?���Oc�9��Y��&��p6����[�C�N`�{�Z\N���A��Lv�ĩQ篤��jX�;=��-�9���ugQޚ�>#��4[%V����#(�n���R_=��>�T(7Vp)�3�	�q$Q�?�y�zU5��,����T�pm��d����A3����^4��\
`����Cc݀����21����l�_�\/� mS阴h��@�FHG9�CθV���39T����k(a���:fg4�0*?�kI1sd5h`���RYn�u�ю�^��ְ@�{��Lv��)�j�w�DޠԜ��vĜ^�T�\IP�5_��� ���;%�4��ٟ<���_aV��[�IQQAy��Si�������s٥�~��H���%��p~B�ެ/��4>�}���zpΖP6����iߓ�Qc[�X��D&�b2��[�$G�DfDI�˴��J��?m��p��K)C���	f��8ˈ$�������q�O~*�7�xe��}c ��V(���<����bύ���{��BX�mW!��J�ON��s� �>�k�K�����yH���B�����m�m���o��n��$AsۖD�!痵��k�[LTD���G��:rݭ5 ��P1�K��i�	����WY��h���f��b#s`�u�g��ك���D ��dzG�!���!^Dv@�Y�ll�eO�t! �����3��c}�Ti��s�kv�Qok��mw�՟���i ������Q�v]3����5Ӌ ���ؽnx<��3�pb���kR|�&ru�TX�O<�O��3=ܦ�)=c�� �P���	�k�X6����$��K|v˛