XlxV38EB    133e     4ee{�æ$�ճ�Ɋ=�"
f&r�S��3<��ϔPÖ�Opv5\#�ch{����r�E�q�0��q�(4V�~#]jA�C��b��J'�%���ޡ8 =,�$�X�X�t��%`�5	��z�6�#h>��P�o�Z��>� �W���NkE{�O$�c�A:��`!��I8����~ûb���FıT*�wI_b��ʋ�l��K���8�D7��g�5��Ј' %K=1<�eE� �f^�Ґ�;�$�TEV@K�ٛ��]Gi�uz`�tZx�_�2̬�*�HP�[��ن&^	>�x<K��YR�@�P?�k�;F����`"�8{���;x{��#�q��=���IҚ��sbke+��˝'�4AB0-�Y�8$ ��������.�t�G�O�6�RNJܞR�X�b0ko7�����Tn���6���RQ2q�;�C���@���+*;RW;	�@��θ$��o�t�[�wϥ2jP��	+����Y���'.�lv��t�i��YZ��0�E�ǒ�sj]%5��L�eN=a3� ��.���w7=���^u���ȡ����*���e�vʬ�:8f�@�A�\R�8�3$k��dr���]%�6�w5��rH��4	4Qcno%g�΂ew��[���GՆMt)Cs�6��\�&�9]��s�y�5�a��b�uS���p	 J��ߒ�O��D���
�OqQ��l�2\wT�7;��;�Z0��(7�V ���Q�\��Z�q��q�O~��5���X���z7�5;`N"/:�M���tG��\�����������6u��ڶ�#m8k��.��00���J�@s�^热f�O��@������vWNؗտ�����(3����f~�^�W��ń�
��8V�������槾G��و��ϫ9�`ܯ1a�4$t�_rξ�R��vDFV?vس��rZ�I׼�z<Ib�/V0�WA��i�� ��3�Sj�܆n����&�ן�����
!�6��ߓ4�)����P��B��\�)M��#��)�U��r�J�*��Y�|�+ë1�g3�{�AJR0���4H[�i����0W>���C�<xn�3c�_7�4�[�7[�X�+�?�(�`�u�`u���C#~�I\	Au�G�'�x��p���W�h���u�o¦#�d.ο�(�q�#�����+u��`[���3	si3�����=L}8��2��ΐ�=�'~7]�c�����