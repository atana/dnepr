XlxV38EB    1dd7     649|��Di����<�w���E�+`��n,��[Mv|i2t���q)ƙ�:_���x����6ɲ¬<��,7w�<�k�Uu�j��'k��lyڀ�����=��(��3�;�����y��H�D����Z�=����p=C����f���_s�Dc0�Q�	Ƥl��\�(�r]��%��j�g��k����+@���4Ʋ��m�5���5 t���`�ŝ�Ϗ�$Yy�0��,>|\4Pp��.]�l淿�`v�GΉ�� ��'��He9��X��SX�E��������Sλd8�B'WF�ZF�<�2��hI��K���>��nV׫�}�C+�X���uY���t�����*p�qc#T��oG�	��;�IF�kR�+���	����:qu�@���Er̊�N�a$�I�̊���RH�M�t,�F�?�":j>J�o�##��П9n��X�[�J+���c����f�Mc�Ĺ�3�^�3ݶ0WU�Ԙk���^s��}�o��3-D
�#��!�YP�4b�Q��0!\>������˲��G�Y��T���k>�qy�4>�e����Vc�U�%3C�w�C^"T�7��;���npCl�N���tVr�!2�uТĻ�*�?�	l��>�Ɛ��B�Y��h�U��!T�.l��@��}!>!�#�1X-J4��뽚3^���8-�$Zj*o�4�
�b�o���\c��s�r:E���P�� �˓^!�l�����%(��6�3��(�P��C� ����®�j�t�[Ӥ<��ˍ�h���_��Ԑd��sH��!�I���pxc"	#;p�����*��7�"��:!����v��h�^���O���;Pc�^���zѤT�\q,���)B>r�q�w>=M;G���ԑ��Y)�v���� �^.���� ?ȑ���A��A��;��X�\����:Lչ��*	ct灩0�|S�y=���c�'�ޢ�����C�e���5�f��:�+�.T���W�|����s�������4�T��IC�xy@�L�Z~�|a�0�� ������|���9~�b�U5>vk�H>���V��N�>�U[�e�"��8�z��#��K7��E�*㖎}]5�<	a�.KAeP�:�0[���r:�\h���<�.�{
=30���3�Sr�!�x�$�8�W�Ȃ���>{PIro}U�d4K���vzrF{8~�]Tܙ|����_:�B�����=w3�Zr�0�s�燆k����>�eF�˴&"�����p`>>_Ihvh�e��b�b�<�\_��Uh�w�.(Ză�*=�A���wI�u�.8H�k�B�rG��j%/�j��c�t�0�F3	�9oZ���N����֡��Ϲv���'u!��>�{ ����I�d @3à�>�K����xC����������
�QA�P� �9L�D��Eww���[�3���U ����Pk&��םk�����^��U�V9��E����ԧy
sǱi�R�"������¼٨3/Ԇ�
��"N}zOh
��@���!��`a5a�z��o͙|��˩�?}^{&Cm�A���d�K�c{(�̖{�w�Qz��,by�<����y