XlxV38EB    1e68     674J��Jb�ܦ��&���s���B��L����!����^����hf�-r%�T�C=�7�biQչ�o9��fg6�5��Щ�h��hg?E�c�P�]}����Gz�CVJ��5)X�4�z�S�:��c�"[���RÝ������82|�q���N�R������l�W�v�D.G���q(�F�"���2�1��[��p�l���3F'IR�� %_C�{s�v�n":��s@}�4횜��Ȱ����fǵ]sy�N���gH4t]ş��*!�Jx��Y��Q�T�6�=��vF���䈁
�P���?���j�O�u���c�EN��ܦ��EjlI_a�"8b�◨�iìT�*θ7J`�q)�Zi�*E�y�0SRtqv5�=43�d��\CM"�Ä��!��ed�U�P$R���k�h�:xޥ΢q�z0"��蕾 �:NKr`�6r	"۾150����τ�#%�8l�{RC�[Y���"��}����K�����8o	���N���9���|�v��=ɹ����IRvE��c�_Z�GM&��%�"Hh�+�$�n+��}n?�W��q�S& 6�������v��g������ga�B�]D�J
�)`U��ׅW��f	��JM���ʽ&x�є��Z��˨����۴�３+P�$�X�g���p���ԉ[�YiY�x�S�#Og�"e�_�R)]d�x�!T�ɰ���ݑ.0�Cm�xC��Ζ6�$#o���As^5�`�DW���ex���6�o*ǤH���j��}I3�f���-Y5>����f~�lPp�@l�����YF��A`e��v)0@I�ޢJ�ɀ48�/��p���@ed͌o𗏌��Z'>|�tJT��s�JȦ����cKoK;��B�w3�9~��%9M�����Z����\���4����8$����	�YG�zl��6��Û�[X���Ҩ��%�A��fN�]Ő�u;��nD@�N�P6�8��,�M�D�!���{z}��6�Xih	�d R��1����mfa���Y�~d�}�ׂ��R ��)��1��\���}����B�v�T|��)��ɽ���LݓTa�Й��C���~1`@��/t9�۰�K�2~Y������Y���]XiP�H�B�V2��Ǿ-ˏ���"�P���zK��ӥh5�0�T����8_���ipT/G1�v!WO�Y�sϛ��Ym/;��Ǔo�B�7�Ch$ Gl�qP��P%��1�3 .Q#g�o@���,�\�n f�#K�U�|D[Bs��D�l�9����2f��jIˠ�;�D8V�. G�#�rLg8�[Z�,�÷j�v@҉�G��ϙi���w(��'�p��׍q��m�7� #-bҚ{���U@oɘ�\�g���Re�^iG���c0a�� ��P �$<�\$~��B�!�zЙ��`Ǵ�������1so�Яw�kS����hqs��QS�������Ӎ(����b�@��6�,I;�M]��x7e�u[1�ߵ�K��T��<A������6�VD�=�tK�V���=��̅3�eW�����P�E��n����'��������i�:�ހC�(/�������n�/��xtq�E-�����J�!� av�����9^8�d,�8��I�