XlxV38EB    238b     721Mb#*8s<'�\W�!��6��%xfoX��tN]yu%��=<$h���m�����,;E�hS'�!	ѨVV��>i���iB7�E�����I�����B�{����&��sPr>d�H�ġ�̆�۽�z ��R��I�2Ka�yoPs�:Qd`�^y�\��L�煝d��	��Z���2+A������N%���?~�cC��aϡi����ha`�%C�^˶�d�G�+�,�s_��d��}{� �hF�J���y�'{h~���)�ƾ���-�!|���s��b.F�h7X��ȺvC�uoWʅ�jd� 2�~h�F�N<�51�K�;��M��#5��v8��� |����J�j�&�]kSl�Y�Ȋ"��f�a���8�M2����r�d� mW��<-G�[1+	���g^؞�6EA`�.� A'
�7p?}�"t���M����B��M�,�U�w����>�"G���"�6վiR�Lt:gZN�YI�آ^�T#PDl��A��5�����Z��ț����ͰܰZQjxc�!i���
��ԣ&卅�g-�B�S��!QZ��t���{���|��'*%��kU�Ed�<\�GK��(�?�F����T�	V' tH Z�'�[����uKT�o�S?�.���Y8i��&��!���:�vܞ�� 
�e�J5Kt�sZ�vܑ1wJ�'}�C�\�	k�M������ ?����099W��:����yhW �5�}`����=9f�zQ�fU|B���]�D%8(�0�sGQ��gʀ߭V'��)C��p���P���x�\D/���-f�A�Li����`u<����1)2u�XQ~Q�<,����.`?m4	��^>:�ϳ��v�HGB7,LiGz�����;�t>�U`#�&��0�y��B�m��,�Օ���̡u�K�EC�2���(CZ�.�]	e9`��>
x����K�ޛ�l��Ir�cZ���_pۧ9|�l�K���I�`��E~
?��ܭi��f[�~��h
��B8�%L��{�O�����dm��(?y#� Ȣ�� y��HAI�`&6'Wj��L���7�/�&�p������ �ۅ@~�s/���OF��ƣ��\,,A�7�Ly�TE�	��+���OA��c�}�*��./R�x��l�~n!����~�5>(�Uޯ�~�IR��A8���o%�l>�Ȯ��p����o��&�u�nϏ�I��Ljm~U�3�.>�X�Ii���
������rY�eN�O<v��pk�^M��!�$�@�fM�^����9)�"��?�l�`1������k���Ns���ގ��3��1}���M�G��eq�����ft����F��1S�0 �~��s��p��}�_�H��3t�߾ԃGsX���Ɯ����
��;�U��� q���u3h!�7��H�U���6�M45���}�g�g-h|�	Gk󽱮l�����kr��)n���� T��;v���`�T��T�+�e�K9�M���?�i�B���\�ئք�lF����x�M����F��>j,������zx����3�k��-�/2TK�#�x#b� 	 �y���@��-&��[��&�\�G�L+�վ\j/�cOQUh����������fh�B��<��r�z��(�ߩ9��C��Fe[�����l�?j�U�j��b�$Vȧ۝-�j��}��I^x�"X�u��
fw�=��bU��oς7^y�|�a�����ᦗ0���9��A�0�[e����Q��Jn! �2