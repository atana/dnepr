XlxV38EB    1c6c     700�y8�	�(�X	��"����dk1��H���A�U�oꖳ�u��UwR�P�D�ľ����h�FE��*� �OA�H�n��C���,�ћCK�m�in��41겅�Џ��8�嗧N���/o[Hkx��
�[�߻���a!���tPk�B�»�85��j�*�Ѭ�)�+c~��tB d�ػ/����h��|�@d ��H��`�r�gZO��W��#�}����u���8vĊ���A���z����؁A����ߺ���5���O�~�rT@���.�B�s�^;��ψ�5X�E�km�ð=ܝ@��	�N��ތ�d5��i��\�3�׸�sG3�"C�+�R�	�!"� ]�5�r�E������X8��5}�l��'��#����������|J_t���e�G�B��碔�VP@����b��9J�����<4+���~z�2��
��ս~�j��F�TQ��	S�M�!Đ�t�`W��M����Qۻ��%g7�>�%�u�����H�p�]�kj�L��3>A�"��觹[�|��)/�,���W����0֊��B�^�D
2".s���۰��58a
��X(u_!*4v���δ����8I��1�T%DHi���r�,���£�Y����m<��=-�։K����bz6��o.{&Hd�.d<�4P³f#m��|���fi���Y�S#7~��!E�.pwM"�R��b7���Cńm�|�:;�[s�~&�Z�?sm�`H:/���y��=x���ÆUwk����[�-���:;x��0���SWln *v��u�<�<�[C^u�f�5� ����N?T0�6����4���~t9��1��A�&� efƔ�(�?��Gv����b���KeU�V��Wj�6��=�F�L�/������˸�z5��YCVc߿Z�:�td.�B��@)�;�3�pSp��>$9�1Nh
v,Η%8�w�s��e�$�Hj|{���|v^e��g`'�\�^� ���Qp���l@��\�3)�@�v,e��0tUuF&��d�(��D���t�O���{���ǉ1|��Z��x�|&x��ǭx����k'�W�(�.%Jl�*�O�X�;uNk��>輚�;]ɼ�� ����)�Σ�q������!���PE��+-��I!K��u�R�^*��`/����V鞆T��!�>�`����Ty&F��*,k�V��\;���]�HC���,��T@_�ܻ�D+�"ڃ�Ƨ��Z�J��~?�ޑc�b�#�21חд2��j-����hB
/���R`��)�4C��x���um"pM޸���^�k)��$%��h?��������ٹG�?-N7����:��L��z��^���^l 1`Z'��f3(~o(Ǹ��J�J�?wۼ�d'\��@a����<ˢ+��Pe�s� ���)U�S+��y�9�{��T=9��SԚz�(z��4�QT>҈�BzLq��2XCOG�M}s��Ss��\_(�ag�e�r��Д�L�5G;jW��(�l
W9�'��{O�
�*/�1�_y{��!�Y����0���^���e�#��p�^h��~<����3��Т���l�� ��X�
U������}��-]��y��zd<�W��o�Fn935A�[	R��u���O�4��m�$m�b��69�k�; B��r�_j�~.Q�b�.�`�}��ȟ����&�����X��8�w��b�l��K�~PK�h�����x/#��W�U|Y��5�N�})�k�V��