XlxV38EB    228a     849;���~Q@Aљ:��Cn~,����x�G+~���'��4�<�)��Iȳ&%fC�t��u�G���)��j�����{��3��k3oݴJ:�VR��k�a]$����#IzQww�}v�i�;����^A�Μ�~{Lo����mR���<ע��Q.ܭ�x�+΅騗��9H��zؐ����$O^�9r�sX�=("b�];i��R����!=�%T-��L���_�Ak�T���z����B��i�9�ZY�C�eu�� �Q�_�i9�@�,E�D@��Qk�T@.x�h��ϴ���r����|p>�{{�A�\�э�]��].e��%.�ȈK���xLn����~J�<���1�<�R۽Yeǵuo �U����	�O��C�kǍަ	�>~�v���Ip$Ȓ��R�&w�9�P5�TS�|�)(�Y=�W�=�".�d� �>o&�B���!-=D i(��چ�~����w�U��ECAj�֤q�Q��fpq����|䏷�Iɮ��x�2$Y�s�_��;��B���z�C��-�
}p8�C�'�d�%
u�lC�H��#"�E^�wV2� i�G�\��rI��>��k,,��N���FN�b�}��\ʲ/���~����z������M��Xɓ��u�8:��z�A1S3�����+���h[	��1�N��>�)K)1U��%f8�V�(���j$T��S�����.% ��nS�$����C��/��zd^ji�.��{�	6���e`�K��&�bSԙ5f>�Lޙw����n5{�� �q�[��S6Aa_��t��Khg]��ͲC3zj���@8I7]���ܮ�Ֆݬ�>����O`����|�ɟ�&e�ueP+�l�d�=�5�ڙ����z��Ol�����<���"����Қ��<��-72;is��FK��W��'�x�/�XwH{��f<��/�ysU��$�_�Hd�`9��X׽ԍq:{nS��յo	x���z�����rC]���k�0��I�ŻW�B~0w7���~3nh���;�懗|��5*��h���������� �+c7C/I�P}�m�nh�ec���$3��E���`݃BʜuG2I�c��̢�j������3�=J�D+�kW~�?Mf(f4�V|0$,��	awcy_� t� 3��t!��qR��"m?K2�:֯�N��޾��0�Y�2Y�6��[I��G�H��.��EjUA,�a'�P/�i�_箰c�OB[��p��Tb,EC�M�<��	)H��B@.��e��s-h������4vE2^Mf5L�(ȃ�����I�}�<Ɏ\��*M���.Gi�KK�T{_���~��£� ߖqΉ6I
d�n�_�<��ɝ�p�>�ڸj��c쯐rg��}H���]T��up5U�$��p��օhɱ�4D�����T��$�i�>��ͅ�,�N`�!vff����2rq���k�:��R�����Q�8�L���L��-
<�ʸI嵩R��kT1����q��j��c�FK*0Mx�<M綿�!CWG�S�3F�}�?g�C�FÔyp��G�3t��?�+9�e����}=��~�G㓄� U�(��[$�nr��NǑ?��g֚T����'!�Ӯ�$Z�����`�� ���"Zo=���󸸲��B��0��<��� 31bH��yr#>D�q<検��J����Zz�|@&XJ�Bg�#���3�{�-\t��#��<��?g��isux�Z�	�679�W�v��b���KG�T�����S��4�]��N�z�>-��e��$]�A`��gE?��M3���u�����W�=����.d�j��%h���w,���K����e\yB=�~����Cj���M=�������"_��8��
`��%�Y8�ޕz��} � ���6ni�i����e�X���u�˂|��5�Ż������½�L��G��m0k����w�=7Ք�T� W��~+�R(`8x-{?��\�Eg)����O�c����Q'܂�or���ĐG�:%������E7:�t�����h����5%� 