XlxV38EB    b275    1f9c
�j��a�=p��n���]�uN�k:wr+-Z����H1(�И��$|�^��C�{#�aS���:{`>��0�vL�Mj�P��;h)�Q7#<�A��.�'D^�+���<����RHz��G63�"�}�>Tr��5-�Մ���Q"	{�w�R��x:~�X���j�
��V9���G��4���AO-W���މk�z��Й�� �#���r0�bt��z��}/�n����˴��0��Ӓm`&U$^���`mY���Z8����J~9��E��h�>H�PG�1�ݿ7Z,S+��P��d\�vyS%��)£0b_�@�n��`�������+�yz��+K]���9����'V�
9�/�7��j�+��o��k�����j��`B����`���*�Vj�x?ޯ����a�?�&����/�+6��l���I��_AN��}#V���=�:*��V���1w��]��a6z�{:C�0A���y�_9:�D��.��� ����%2:N���X�Ҧ��~�M=��j�7�F\M���3
ע1�IP�Y�1'�^�ì�G/$dI����`�xJH}��������AfSV�dM�h�G7y%��=� �\�F�b���^���2���" =9�~8�`U�Z�CХ�b�5��K�m�ʱv�)��j��#����T�4�n$���n��� 7���9gG�,�W	XrIk��Y��Dq$S0���'X��8��1�<���?&f- O�P�唘��켙YE��LD]���X��~~�]���9�A�^!���Al՘%����$����ԫ�xP_�Q��#��/�<[���7N��[`��~�-�f��p��?�^ǹ��+J}�O�,��7���c����]��\iy^�d9�sr@���� ����s�˒\޽UQ�^���G�ʜ����`�]�P��Y�s�E^�K���	�a�]��yG�ih�]]�@��-��jn��c�\��5-�EA?��[�F�qN�dS8×
g௴�����Kg��l T�O��4MQ��FD ��G�Q� j����� Mʪ�Ѵ�;9֧GtSR4�C�pD��e�X�xd5m݄��):Q(O�`�=�~�����1��o�k77
劀�����I����~��_z�'ރ�@��>۾'��}8��NP��u���3�͜��� 5ͳ��i �d���B�?c`�@W�w�����o��f��<K4�2G����j�$t
�6	�t�0�ǻF�A�f03���>�#��q�]"'�޺�|���L�7Ex���Y�R��o�6Ti��#j�N�r+����u�K�6tQB��-�Ǟ�}�זm9'&�_*J�q�k/�.rW�
I{�C[��`�
��r�2>vpԌ���qolжl�H�NS$�qt�?���*o���Sq��m��M4�S��H�&9�!�o#7��C�)��-E%^�/� ,�Ԏ�53o!��#7�<��О�fbk50�҈(���s�G��)�s`pz>sӢk\g~DA�G�i����MER��.���U�yǹGo,^�����NE��[o�S

T$�c�h�'�����49Z�Rp����fۋ�U(���z2��T�]��y��g똖?#�p�UB|À4��U�hj��Mm
����\�O����d�5�I;#1�@myYc�F������h�w���mj�壐����H� �����v~��_|ԭ��$l�?[���V}�S3澢N�wVb��u�:coJ%�$z�����%T�\�Z�_m
T����3��>����jT���ς6�4B���E���Q�|��v�,ߜ����]����̰R��Za�#e�Y]|(����7�?���r�v��$����͚���W�#�xs����D\��U��c�'�ڪ�p�`�@C���7S	(H���vq9c�e�W�+V(��aI�x�0����=�oR;|����m	K@�Dk��x�$?ϤX}8�IL��	�ܙ*~��Ƒ���,ď�����<�'?��oT|��e><h�M�C���R]?4��
��<n��D�Z1V��[ns�_J��I�.�����T�H\5���fc�3;����7ŒZ��Wqm[�>������ř�|W�&�����9�o�)B�~]0.:-�:�w/����K��ڌ;	&Z�?��֤E�t�Y���S�����qRҮ���Z��4W����>-!��T�̀02���9~��b���o=&"�3�/p�B�q�v�������Z[U����Mv���h��f����F�&%ъ��D��ȶ��E"5����R\-8JC;n���WJ����G8PМ�@or�rH5��,")?2I�?$�-��O3T�j��+E�s��{��Ѫ�i>/�ś咉�G0T�*�ːkl{�Koj���	���5|g<O�5��A�'����-�����.��x�7)���2%�q��K�}�/��gw)-�w���:��\CO�v����.��Q��p�Vz��&3Y,|���y�!	T��@�gK0��\��KE��5M�	��!.�0�Q԰�K�a���&��U���Z�;���?�8P���v8~����c�B~��T�<0��I^�,G:^'Mh!��i;�f/�W-�V"0A_.����*)X�0�������ufO�t��R�7��/R�(�^�K+v��,LtlNHv�>�o����$�Cb`��w���+�s�Z��2�i,���h�哫�����4`�^�	��To��G��7�`E%�`�LNt���(솄�US?�q�R:�G��\���4l��J]�K���l�ЍA��5.Y�h���ߩ�2!g�z��� ��z���"���8+��7h�;]�	�(N�S���O���Z��:�����_�R��l"u�h�y��p�߼׀����L�yT��,�%�a����������I_�V���P���`��I��5�~�k�)�LU��;��+�0%k�t�YnB��}�_����颸���/9��w)GS��7�}͈�'��B��5V��72t c�ϙY�������b����E�qy��
����R܉AAR"@_�%o,ɜ�����Cns�H��1f9)�j�ZG��g�'�c؟�,;ͯ��i���C��:�h㊵�5'�x���c"̣Q�F��4�*~�n�}��>�2���'�	MB쇧μo�EQ*��n4�L/@|��q��&��"O?p��rC��!�	*!��dMg���<����>W����ݎ-B6`�xo�:ݬ�27\�޳}�V�`�O��N`����1�e�?�=J@�����c�r���� ߳�zw�1Y��*���)��u���b��v��S1��wׇ�,��fl���2�,0'sc܁� X�x� M��g-{6��t&]3)]��AnQ�����ō,)tMLC&�
�����U���#�8CW\ݣ�rJ���K��3).�Ҏ��W�B�[@2�
1��q�������0�ܹ�?�[��ޟ�M�Y�p��IK��[Pϧ�y�E�l�a��ng�!�v�K���輬����fd^偊nC~e�՘)���;���gBBȬ�����uD�m��B�~���}�'s �"iBd`?�G��XvMU�Qp;,	�0RG��5�}a(��2"�y�+)�6���A�{�S��Ǖ�,�J��e�km �K�.����^�,��@w�F%@7a���g|�"�h�����X �mS��W-c�j��o�ѱ�E&M@V=�`�Naw����NCTpQ$x�L�Ǘ�Qw�g.�p�b�Z_������MX���~A��'?H��IQ�/��{���|�6=��.�������yG�l���r8��^M��ڝ v��*'����M��4�<��7F�����X1���7v*>�8�+	��|UBB.�i���	k���5"O+������|H~�ޚ(S��O��.hb�y2#���{@������Il���c��n���M(q�#?���gQ�Ȉ��̲΋ ���.x��Hr�ȃ�=v�E��m.�ήA1�H3I�
�����"e<Bo�R�:�䨁�5Wr����YS�������uu�%���sU'���N`s�u�>�6��|w���#1���S��Z�oG�C|��iV��_�����;��0T$�����7�7e��Jp�}gϦD�F�rG��C��9��i��� Gn�7^o*/-6��	=�U�s �c�C���8�PP�m�y ��03�c�a$������Xߗ2K�t�Z�z����j���l�`q�*w�_6
|e=Hڌ�'e�m$�+q�2\���{��{��i.%��>Ԟ�g$��Coh)�� +k�@l���%����\�bS�Q�l�_��E���d��)�G�N'ų������i?z*��9܂�ZA�}ڇ���^�z�HP��b�[�[R50��/���s{8j�X<=J-L��w��|b�(��V�އP��Ʀr� F��CLC�.�{��9�)
"�FFIx�[��	F�}[`;P+ ����H���h����%>jK��}%��cH"ێ �d�;�b��7�� <�"7C:;�cX�}���SZ��G'6��WFE�K��f4T��	6�����hĐ_�0�����=���<j�����.�;�I<��ȳeګ5Myf Fg����?"�
U���1�C�}V}ӆ)<*/6۠?0�mva��z�� �Y�	o�l��:]ZEJ�3�-�es��e�"�]��1D���
p������@��=����7����W�6"���֤�!ă��Kۑ�'h� ^�N���>T[�ט��4��Nn��G܃�ʕ�C�I7F��xB�|��Q��;�cwe"Cbp~����q6���Ub���)զ�fn�v_S��!�߀��f���w�km�ɘ�E��k����P�)MiY�_"g��9�U�Z���;�<�`*�4���
	�6�Z�i
�yMP�m}8=BCNN8#��<4�}y/���'��z��K:�	G��5�U �섖�椰�⺕���kOO���@=�[k�r6]�n��%����D� �/Z��Ȃ|�1����M� P����TU�1Nx5�-������,�.MC���> `Ϗ�J����>��\�k{�z��r�]&lKЋ��� ��Mg2����\�	�H�t���J �k xG���f��j��k�$52lS����$<��{�x���x�n�q>~���p�(��vYl��sv)�m���3�}HG�aa�J�^�9,����d��TF���*ت� ��7ݙ�����o��͒�"�kl(������ΐ�-_N�@M��IeW���4!z�ҵ�L�ĩc5�F������� ��� n[����a����g�ʍS*�F<�h|3Cw)�5Fi��P!��J��� ��B�#Y��ǖ2|���ŕ�����Qz?5!��ݿ"�q�`7��,�J�>�4�*Z�ox%�H;���F���ٴ��a���):����[.��)�O(�d�7�n�a������e���d�3��/����h�zׂ�M�'���ejf�T�4�v^�%d�Z�W�㲿�9�[Loyи�~�}����C�\����(��PX4�/X#H��8�]�wk��d������z�(j>�)��3�d��f��������W��>S���BW�9V�2�o����F�x�ٓa�Y�,��YQk`Ɋ����(܄�z���B![v�4+;ʘX�s�os�wU])X��Х)J�ǉ.h�Lsq��	�v�r�d! *�;�Q���uw�&�vM8%K�r�	��[���A��0�܍���ܦ~�a	4���i� .�,\QB���b�U�f ��~�Ȓ�Ͷ�E#��i����N��"�D�X!Y.8D��w{����%����9	�k���ݔ̂t����ԫ�{�S��8�S� ��$�R"i��K�1��bm*�l ��|cT�tuD����7���I���#����=o��������o������D�w��dq�)O�����������S[�%�w*&�6��s�F�J<3^�+M3��4j}Z��1���w~=&#�+�i�5N���1!������|����`JU��Co���P��>���S�;��c�c�$횗V� ��;�����R-�Xb���?� ^���[woTG��|����)Xs��<Ut���jAj9�@���0rp���S,�U��#�*8G"��p2P���73�&KY��.��[�PZ��I�!�;5�<+3)PQ�9�/�|q�Y��$�=�Zm�3���m��gz���${�vN�W�:R.�[:#��%p:����?�.P(-2��(%��_jj�Z?R�~�;��mV���P̰?����G���܍ֹz|������ƲvT:����K�m�QPX�7}4�*��sO�pj���V����Iĵ״�-�����,V������;�L�R�l�yh���bƶE$��h���?`�ǃf�1�W0�+2_g?"��Rr����d.q�_T�(�bkC���\�zPz*�ډx��5w8��A�6n^n�+�_1Rs�Y�EXdu$Ôp�Cq��|��2s�l
]n��F�(��+���Λc�m$]>ٺ�Ƶ�f7�+O>"^��@�?ؖ�j��]D��ٽ��ނQɤɇ�b�T~�pԙ*�f���pV�AAĂ0���|��Q�d�_�k��I�T�����|$��A�	�����+�1*�}��f��k��+�������ֻ����67U��$��oL����@MD��uT����{�
Cp�HW(�)p	������G�]�jUj���#ǉ�q���P�#�������*ۦ�}d&��>|��3�{|!Z?LN����"�\�&��?��}A�;~���).@���âS�T�)�~uf������ �;���qq�¦%�)ى�K�╙]H�˭)
JQ��ڟO������js-�粗�7���]L��d���"?PS[����3*r���pZ��m.y����?i&G,��j��&ގ��k]۠�@���^O���]�.ݴ��C[|��KFU��Gy}�r����Y�BQ��L���|CDג�W���J'o�������HX��,��'/p�0�p���I�U�h�����o����M
K��@JC�`�~��kWT �kȠ��/A��X���=��/<�D���1�O4[W�>�6g�>�-\8x�_��t7s��>{	s�\՘���rݬ䫊fp'm�9�1v�ڍ)U�n�g-��@��2 �L�SC5���!�A�^]/������b�$�$]�������B��V�$!)��f7����Pq�.���g�l��I� �B!�	�H�G�>�B'�a�7�M��um�1N)`6�D��a;\	��6Q-�Uk噫u��_�>��8e=���9Zcl�D�/�m�A�v�W�m=�E���h�\��)݋Ѷ$�*Qg3@�3�Zӎ�f���%~~��ϥemv�����1�A��/,<�Tc�xv�I����t�::������_��RC{n���?Ѯ���(���9�jcj�W@���Y�q��'�c_ڒ�����pk)�{U��[
���u
=
�@����p�y$��?ή9���P'�����(�L/F�;dܪ)i���˜���K~R� j��9.(�$	u,Y�S�(��X�8�O �uYq�:�d�d�(�[���u��"�����[�K��ۋ���pO�}v���~�2�ݜ�ѷ&�0��?��*�22F)�Yk�˃�oG9%NAl4׺mv�~�i<���[���Ȋ�V����_'��SG�oo�����ޔ�i'�6�ʄ�7?�z��Ф���Q��oR���	H�BZ$;�5��ėl�4ݵG���3�-h��>�7��Ԙ�A�.֡e�/{]����K8DK�IG����YӾ�]A�0|