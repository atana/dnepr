XlxV38EB    207e     a2bpW�]��Fu/��?�q݆(R�	��!L��K��������Ƶ)i�pH�>j8WWh��ncљM36µ���1���9ƿ4�-;�s۹֖�<�ҿ. 滑yU�P��?�4�v���Q�P�ŕ�9���,�]Wz�q�R5���F�v\`����g1��_�:�(�3��*��I,Z�"������D,�2�Z�u ��e�*��_s���Z���眪�����o�A�q��<��[��\zz�ߔ,;h������ma�y(u'�1�Wer��L�;9�sC��*������Б��i"\�̂�;s(i�=7���LNbZ���mE�	v�I*n�
v���r`�
�C���WZwYc���cg�k��ɲ"�!uz/��t,�*�?������8e�7���!,C����C�e�b�խ|��Lc�a��.L���d��B�Ĭ,y<AN����e����K���Ѡ#>����j;)e��(Z�JJ>xXQ��"���/Y�0��}�$�T���-��st�h+���+O����������	m��OjGo�S\G�̎Y$��!eI��ZK\��zJ�8y��rT����R�_ـ�i�Y��88���Nnz?�BF�be9�xQ,����Ȅ��r�j����y ݁O���Gy��j]��F�z��|r����n&�4I��T�g��(�8Y�FQ�<嬂[=7�p`�+&U71 'L��j2���w�q�VZ>���?�����D���	,`��Qڒ�P����y�D�f����7G�?H0򃍮��%G��x/4n>[?�eZc`�p~Y��U�֝�\��M�Lv�:�K]�o�xcX
!�qA��d�p]W�{f��W�;ANu w���Qs-Ӂ�@���:��9�&�I�xyƌ�y�y��@��Q;ͷr\�!��v\'�]�rF�i����،�Ѹd���i������v��P�V�f��U_
��@����\<sMfFj� u	�lH�E&��;��J�x$8]7we�pх*噯!�+b�I��W>�}�?�/��'�0���h�˞}��b��Y�*,ڋT������7�����r�[kD]�T��?�n�$t[�=�:m����(&�'cV�e�ɜp�H�*���ܭg�B���?p��f�u6�"c�b�X��ܜ�r%�ùᾼ��IKdپ��e8���!�5������7i��=���D���_�v�3ä�" :.+�K�m�͏i��?���E���bIü��&k��4ȯI���/5ec�W��C9x�f�0�u��Y/�'b@����Mt�3ʷ�B=IE[���Rݤy��;Z�q���i�E��IUyr�?�����n������6�pD�wI)��	.��a{dX��A�?y��9�R]}}���8��)��-�f��f��2�;>������0��q��2P�N�ެ?-p&IZi��eݕ��B^N���J`���<�$0��²���۹�m�&ԞX��]_$j���%a�̘�<�x�= E�v�X��� MB�U�c���[k['��z|ú> �)+w���`4�[����%�$	�����o�����f�鹭4�ח�ݖ��,f��)�)g%"%$۵MF���j����Q �!p���d��sIV�4�/[y�y/%�F�^���ܿ+@M��'����@�J���y�o�U�kT��8Z��E��$�	+H��f�:���w%�އ�t�=^�ZQ=~����?[��ig��(u������k��b5<��$�s��7A�8�����y��W�U�ᕉ��'�\�e��c��m�Ͳ(k�';"jM�xUr���F*G��
�NHiR�:T�2'�OP`A���g��i �%��CT�q1����1~r?�^�C�蓋�9�l�&W���Q����������ho"P�i�~GO�#$I���%V��s\�X��h�n�buc
����4�n������6� �w�
��T���d2$j��&�0�ܢ-�3�W8��j+�q�4,{>��$��Ȋ�.�I�� D_�r'��#�P��nJC~z�q0|3�������u�j���͹����"AM&	�4V��b�
�������mDK�	�{�{v$����]=���*�}��Zu��d6�M���g$�W���MIO	�$߄p(��å�B��Z����7��������'f�)6�m
��al���?+I)���$�T}(�Y Q������}Fs��E�՘l,ɒ�+,d�b��E�7�ƙ=�A�-J�w��?��r�篜*���s�@A�Ш����E�����	UI  q2��<ʮNX)�K^ç�i�R"�uJ�[u���Mϸ��Fx������}�_�uk<�*��̢��/�DԀ��
e����Zn&-	����x��({}�x�f��FF�����jN�w��3�vi��B��GG	��d`C��%CG���Ռ����ܷz�qE* �:D�<��o&�&pr��6�	��1��K�P�s�5���aƢ�V��ǅ��m��f��^ ��'�l����-�̄�V*�0S�O���O!Ss��SN��`U