XlxV38EB    27c1     9d6ڠ�q'I�3,��6��+��!�����'��7�\�4)�q��lH}��y��Un��x�����lW�a��_I�xH����+�Q��ȟ���'Sl�0���Gԩ�Zй�����Y%t#H5���Jd<k�R�19)k��� 
$aF#�C�N�>��D[sm�I��F��T޽��m�L��ҵ8%��}Ø�����L���2G����[�����V���Vź=�:�R��!�%��L_h�����1����!م��j0�ӈBl�E  �����[��ݟ\m�����8�`�E�3x��˗�o�㝏·�����N{LP�[���P����ڴ����C^�aY��P\0UL/-�y��_jC�+�,�_����<7}���Ѷ�䈧����7Y-�e�ڽ��wx�w��u�2h7�h��`���/��Z�35�d4�3���"�!�̯�O��\f���5=+\#^���s�%��6��u�-S�~��PC�/1J�'d�A:����{ɋ�2j���T��a��a��Y����t�5��Xn��������aF9�����&&,�{R�� ��@��)[�j�WC�x&�XZ�ԉ���]�*�;�Wf��O�k�?��p+�Z�m�uЃ�^t�E/%���J_=��8zeL'�ѳS��	�o����I|Oi����f��}>i�X<N6�6b�z7�~��f�V-7���: |1ӷB���n���G�%0��/�%L}����;97GZ�R��ջ�N*�o��;�e��m
�k�g�@`�:�~}�9�����"��=��a��hP����`�V`_aJ���Y����LM�T^��)HT��������XY9�|������ו�'�4��D|�ӣ=��35tٖm�?j�-���n��yW�ǨNn��<#d�E�ϕ�d�"����h�lH� 9�j�� B,{�<�6�ȓ�^,�39�C���X����P�1R�1Fʮ������)����������1�y�$���QCc�c �S�&A�s���)�ѿܠ��Q���sK5&�"d���>��s|~s�]A?4J�$N+��.�uuo����q�U���6�Lj.���)�k]dT��1���#ͻEq?;N��z:��׷����4���_���+¬� �(G��A�x�w*y��o6G~J:G=�<��-�LS�S����cb/bf�ڎ��P�Ӵ���@({��3��_E҉5�;��J|��n�f���=ğp-�^����+
i�3 ���\�2]1���-gU�q>p1��\��l;�?��Y��z,��G޶@Px�*-�����F|g|���&�{��Y��;�;GU=���٥U���8�D��Ј������E%H���JH�-4��j�;k|v'��3������-:ћ7�j�=p^+��D�ާڎ���4��uq87k���P�[�/�@�Y����K�k�����}
a��"]�-nN�!TK'R��ra޳V�ƆǱ��)JI����W^�䔗"z�W�[���Cg�����"�<<��w8�^�4�2����(��	I�뺃��@�HhׅS�
lPt�1��I��&M�(�feE�8�k����W��P�P8E`Z&��D^�G����Vl��`;��(?��&�9a�1M��tp�	�igfd[�Cب���M5B�o�COt�	>�������y%u1����_P�<���J���¶���A.悧����UqZT�?	l	ˋ >�$���+QȽ"9��T�&0���ְg��̡�&��9�{H��^��q��&O"�u~�jX��-���>�]:�����.�*n�CV���F��G>H���}'|�C�bQjg���9��t	d����\��
��^�0 %pГ��έ�����������_G9�|���=}<�P�����H��3�(#�׉����4�����gk{@OHe��6.T&�F�촆O�o&6~������Sѭ(�L%?���ZB!�Lضsu	��%TCM��⺻�J0t����j.7Ug���d�Y�Iv@�C���<Ψ�"{p���̏U����ȁ�7%W�;L�3�W�|y*խQKT�,|�F��(i�T'W�1��,��@m�[ڔeP��������Rϊ]����6c8�� E�cf �/@�T�.�,y�y��~��2k�p���\?m��q�-i�c�w���ƾ�a�pZ�h�O�~�ſ�:���f �8~�%Rf$�K)�"�~r��
��L��잱��|��gn#�0ͭ"�L�8�W�	�˸q�aEc�'� �����DNO�È#�`��W	݆���X�pe���^ Z�ZFJ��iP� 5�K%q�SF���i
H��ة�ۺ�>�_��E�EF���u+��z��RAbp��ķ���O/^��{;��Xu��r/c�F��d
����M������H��*BeU��6�<D��j:2�շ