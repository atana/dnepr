XlxV38EB    1ca2     658E�<�'��\��Wr\�x%����^Җ>�k>K�_= �>����	0 �72�YI��I��7�H�k��>�u��d�|����z���H�|AS��ZUX��Rӛ�OM�A���S�����I�����Z�q�ɩ�ei���@_ '�C�<�Α%?�A~�n��&��P��ć��,��/%B�a��Bx�}1AcM6�JsgKyp8��J	�J��]{��?V��#����u۰�d����}0WK�|��Uy�L��iiH��&{Xy�F�V�:Xpk�����K��	Vi���(�2�b75��"��lb�q�v�`���6c[�6.GhT�ǰ���WX�Rxہ�O�V�&V64������2���kZ���sA�X^W �0��!�\�Լ`�	�p'kL Ƅ���{�M�m�b���p}���O�&��a<�Z����<�ܓ�+-� �{m�M��m`ǲ��s��w��\ܱXWq�@���7k�v�����A\(,vpo}��?���$�Q��'�~�5��[�� �1�� g�C4aA����l��On����m��Hm�@Ƥ0��t�e��Lŋ�c��9;�i;�n�Z�:1xʒ�ı*��v�����aL��Mi�@�6*tk���J�B�n[e�PBs�R5_^�{F����w_��E�Z�b"��WR��XQ�E*s��Rh��̂I�땧����SF& �꿇q��"�
R �%���TΘ���'�4Q��2u���mh��kT
En�
/z�����:W�[j_��7]��������#�O�����z�b!��cXUh��<'w����<	1%@P��|��RƤ���G��`N�WU�!�sՄ�g-ne�P�-g�����N�Z�"x���R,A��iBm*#Պ>`V�O�.�u�1�O�\Y/�L3WR��\�Nq�&��C��2M|z7"�K�~5�!2D�cӚF����2}/f���:K��B�_�<I,1�j0	��K���0x�M�߽)�U��
R�Z����PAG�2u�gBp?j���
�`��bce)xp�b�9"'�4��x���x��<�G��<\��Q�߲"uQ�n��w��!(��_�]��$J#�<��qĆ*�< 0%�ʦ��޶B[��Z�*+i}1nFt���f�7RR�`�W�3�M���j�b8�|NOpB�Uh%�"�Sm��X�*��R$q7̤����e����"WF��+�8�#_�+;7SY�Q~�k��! =������*-�(Jƶ}ya
?������ūrn�f��E�/��3��$���	�<|���	�5[ ��:����MZ����s	h�:i��	5d���[�2D�)��7=���u1S����n�'�竊B�Q�"7���Z�f���:=��y�g����Aj�ǃ"�H�|ls)%��M�o�L����)�.#P&�#&�٭4�i��&3GA��dsk��d�����~J�;	�\N�H��cQ�*Ȼ�z-���F��p�$�����y�.���׫�g�ذ��n_�y?t�e����K]/H^I.��fO�9=��3��x�u��'�ik[d�p�z�hv��s�Y��k�a9��]���V��/�$/�d�ҵŝ