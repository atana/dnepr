XlxV38EB    12d1     4d7{�æ$��h�'��*1���o�w�x��H��oC���PՏ)�������'ϱ��-��S�@v��j�
��*l@kM��8�Ҏ��8g0�����m0�]�b�x� W����~���ڒEt��a�* ����\./�X���kl1���O3p�U��Cէ#r߯z����{*/s`,uL$]��9�wHr�a�!�t.m
�&�k|�2�kw�o"Tj�8�z
.ĭad�����J���چ�q&���k@7��/�*l��m�g���	�{��f�����8V���A���'Sa����tY���L,=	�k�������x�h��'�eJq����<�<����hEe�YJlloㄘ��Kl,RԦJ?�Z<�H�7�"�W����Nynr�xG7!�MX[�7�1�b.����wc�.n��Qʗ( XELM��Լ���ĝ�C�:��8k�]���ۦœc��?:�@���FZO&KV[�~���<���W|�^���r�8Gz|K��7@TӐl5Y')�ު���܍�P��:���,���{+j�5$M��8�g=��#̋���nw	�A�^
�Z|���f���!��Z���y�v��8�uGQ(t���2����T��~��� T}D�" E}��xg����VF0�G㑑'����43��+�Ǣ�c�Ō�i�x��p[�k��?O�	��)?{��҇C����� �ϪH�xp��	X��Am��Q��I�O}�y�~[��4U�a}��w�'�0�����T��VZ)��N�k�=���D03�~)�M�i�?�C����uC�����kA�~mF���r�Ƙ��K�s�c���!����"��AM%G�5�۞v��sme�ML��&��{$�-8�))�P@�Y`�{���A��o@�X�F�q��H���:��^�xY�s���O�v��b�x��@b9�V��y�S��)�U�cJ��>{LWs��w))�K9tNr�E���m��v!s��x����~z4��P�`��򠙛����|f��E������v.Rrs��M�����y��31�A����4��h�#_�}'QE��z�W��~�T��c�Y�J���P������3�5!	��ƌ��cG�U^�tL�e��et��B5V<l--�q`@��K���C�1e%�5�1�{��2E�\-\G�S-���Dz�1΁xc�"
^9�.�W��p��