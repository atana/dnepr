XlxV38EB    21d0     810�mV�����o���Q��tpV�Zz=dn@��/w��<���:Fnq$�$`T!�:��Բ"�
wOs�!�8�C���������5�4[G�O٨��0�/��N�Ǩ�R�$�d��:��{]�C��)�:�5��(GƇa���}�o���rJ`ܽI�����B���}��j�����$!�N �,�hWҒ����Q����lx�':hI���u���YbG+-��fUǪ��g2R���԰׬�(g��ö/�Т^u�en��iQ���N�=J�p7 ���y	��d
R�Q�a�U%�ݏO$��K�׍�f!	���,�_J���|-��˭gp�����ha�(����F�ٟK�˗�����uc�����'F"[�1�ay�	P��yܼ���l0m�s�R`�!��Cd �����:���4�
�V8[. �"N�
9�X}�|eL�s䯌����c�b��wî��������m\���v)W�V� ��3�����~ÑEK�C�0��r+��[�$�qY��Z�i;�2`�OD�B�-�LC��<��,������z9Q	0�D�n"^��"_��U����,AN	�	`{R��P�)�x	>ˍҭ�prS�u�P�D��T���cA-T��Jd�-`Z��݆@<�~���'�+Q4}��4���v5��{��E˛);P����7�'�'�z��o�R4��&y��p�ѣ!ǎ�� �n��z	��Y����~�"�ѯ�䨘��S�6�yB2N���Sv+��X�[�%iT�
�NU�
NK�1��3��:F���k)�I��(��
x��U���ʱ�NH��ϣuSm2��7������]c ����%@���(ϩ��/��%!�?���<��dR�����J'Vy]�P��c�������W�b��{3(�ދ>O\@��źn�����x鉅�FS�$��]�������w�i�d��hX��-l��bD�`�ua	��Z���g��n���B3��Nf��JK�Cd��uv䯍�çuиMTVތ���X��w�����b@�V�3�
uQ��4�+"ѺuEBԌ�:r}LG��1��N��=�ɪ��AN~ݲ��UW���l�@����JÝ&,7�yj$�����w���,`�a�@pKg���G7�����k')7�fi�����|8�@c5&C�����a�j�m���k�3alެ���ӐJ�`��Tx�򫊏]�sRD7'�!�O��_&�.%�fG�#�dK�fՂ�[� T~�ˢ�Cl]]�+��	��[ܼ�)0}碽_��qCt˾:̀:�)(ߢK�;.vC5�D�Bf�e�r7Ǽ�u��7�LO����/��:���23L��覵5�����Ew��:���4$5��e��o���=��&ΐ������!x��'V����`�Ș��ҏZ+��	�D�7+��+�)�f�_���QP�NJ�OJJK{_��L,�QN��i�7��3[y��T5*�u}d��1����6��6I���"��#���1��D�9�4����b`�^�WN��ʳσ�����u�#�b�V�L���Q��D&�?��������폾�P�^�Ѭ�c�f�U㗜|1{�y���q�,�b?+��5�U	uZ�!�r�^����n���qr%�(�9���(}��˺���ЭāE���t�n�#��%J�{�?����o�b]�a(81�}'�>�7���T�y�k�Zl/�g�a�Xi��~�`]�.f��{��N��ۿ�D���iK`y����N�U���O�����@�a�]�:��̌D�S��ʏ��q!H5Pb	,�p����_
)5	/�ZҀ ō�%�_��b0Sv�j�6����d/�7԰��+|�!��I��Z�����.���<⨞�Ш�������9�F�k������|⾘L��]�*��"��Zȕ"�?_�M����l�,/���`Fdi��ޒd� �"��*Q��^ժ�j���cC��ogl�7E�|���2����K�u�<D�����K��