XlxV38EB    1610     553`P,�3�@���R�;����V��m2�#l�����..=i��iY�a¢� gz	��� 7���g9�A'�}���Yyk����=~�cG](���Xʁ(I���H�]�M�8hhq`�)��I�S��.�8�8tIn�@��7Y�t.o�LTwZ%�G�}
6_ӹ�r�>��-J��`��z�&Q���>�w�<�^Z�L<��P�g}B�(��xij���:�z\�E��l$��?�:ϐh�����7H�̹W�(r}K��*�W�=��$�wi�{��Q�q��,�Ĵ�o���Fñ����2}��!���+�g�ݡ�©���˗9FIQ�,<r�*0	�� �Q���@�L|j���4���6e��!-vDQ��j�	D�`�ɑ��u*~�0��j����Ф�7��i*H_f�� ���L���^m�"&p!M�T�qf6{��y�nk�Le%S�nZP�a1���;N<3X���++f�bA�s��M��*�P��#�Rc&��v^{|b�Xgt�N�P|~�ko�U�=�zU��Ɩ��A����k )�����D��߄�{м+қs�����"���]�c�#ez.;qZ8�nE�I2XC��>�:�h^8���P��0� R�kD8���������������a�r9�tp�A������ �˩�Q)��/�\	�h�C0�K-�Q�Ǣ>8QƢ�(���.�ȳ<��Խ���K4������ȹ�6�Җ���}�T(?�S�W����$-��fwp��3DO3�_Z�KJC�u.�����
�"ACZ$[���`
�׾e?��7�Fo����E�)�̶H@���B���˦_�'D��%*B��f)VˏJ�N�WB.��CB(S��F?��[n��H�c&E-~������q�?3T�T'i��!̝!�"%�����/1�^�߄�D���JZ�.���(\�Z�#זT!R�v{�������#�5���lk��Zr�$R�ڝ8�j�%O�on�d�'���Vd��?���Co�O�XO���1�� ʠR�m�t�����Q*��Tf9�(1�N�L0�V7�����32��(��3XGh�߀N ��zc�x�9��F;��36�!����0Q#�G�:��K3g!`�F�ߧ:�����2c�	��ю�������!�S�8��W���ۢ��������	R}�0Lp�9.p�lj�`Jg 	�j��st$)�˳��qt�����ȝ�#��Q7f+�+V��9�[K�Н0�G;&E�5}��Kw�^���R�ǳ����i���q�=�.*^i��."�*�4�,R�&�CI�f����d����ܠ=�����WƈϹB9