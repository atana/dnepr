XlxV38EB    3c73     bc8G�*L#4�{��T�l���,P�"�3�ZI�ك����G�^SnI5����P�I�����m*�W3�>X\�Q1�$�3�A������H �Ͷ�N5���Iu1o3�67�v��&F(�6�Ӟ'+�؊�k&m�9�A�n�b5�e�u����nl�/��*�d�6���f����K����L���f���q
��Ǭw�n�<�󉼼�(��i�v�2�K��]uKc�X�Ak33ӿ��A�����4����K�i7�����,T�@˰�H�=:1Ƿ>C#d����P���1���qs>�dv��wR<&�ܐ��N�^-o"}� .>���Ց�*���t#z�������6�1_O�=׌S��5]�n�E^�Xc#��?���Lo��#����@m	�;c������^���@J; !���%�O��0U�i�`W��7I��&`&G��^X	��s< l��aɚgt��@�V/��=>�T��Z���Q�q��
���<��T1�����S��v��存u��E����%Ae��SnT���A����U��B��R���Q�N�MMS0�M@�}ˌ�K�a�U���-D	jE��}F��!<�C������nE�����UR�g>?��M��tk���pd�y�>��ce��u!��c�yb@��?�XC�� �&C���v ��;����t�(��ҩ|��u{<n�ԕ���;�E�EY1�iԔ�6b%Ɖ������ؔ�(�-�DQ�Pn�SN�	1 �igY��Rl�+t��q�2߭�+>����nm �kOW�ɜo7[��줁�x��Z51�x�;�d�ick����ְ��u��2���Ɲis���8"iK#�to%f}G����V;�o`��n�1jz�*u_���o~Ś�θ���`Dp%���Q�ͧlj����L/I�( ���i�ۓJ�zQٵ�D�	J� ܐ�*��=Y}�{��}�I&Y[FY�6��Q�������������QöԊ(���-S{��淊�K�2�Z<k�K�}����gA0PD��_�-E�^��u�jx4�z��?�8I�ÿg��|Ħ)�_x ��g�o�v�80�>�M٢�]�\w���?��'4-T�04�-p&ɉ�c~f�?���L���ĀS%�s���&�Fdq���=	�Ldv����PQt��f{ʋoN�&�<�H-?U:*��������|�K�s��҄�>H#���47���o��'�$�n�,).75	&�!��PB1��̄i���=6+A�����$B5	3Q�A��r��@Ͱ�Ɣ�*$�(�a������MX�]Q�A���<~p֕=��f?g��"!lG7T����s��8��8 �=
����@�
��,�[�h#��[�.L^=���c F�G�������\/v��QGqo��`J5p�Rj�ң0���mߐ�!�X�gN�II���)�ʑ�����"
�4q��ځ�!�K.�;Hg�$?��y:���}���!��)G��T�������7�Ա���hs�����;������6�rob&�=�Ϳ�dە^���Տ��c��%ψ�XoѴ4"��-�����ujR�l�٫��t���x���c�g��~�h��?����ǋk�\����ꖪg$����Y��8Ԅ���O6�/J������1���1�t̘R*���G�6l�{ �1,��C�6Ns}0�e�i���D�K}���o�
�q��(�ZcL����Z@�W-�u��Õ! O�IT�*]m
��?�+=O>U�a1����'	Y+ѧ�mŭ²����k`ڍ���ȗZ�E������	��lp��Hu����'y�*�x��b��HG/��aXٕ�h��@M�:I�NP��jpZ�_�R�iw�f�$��S�s��^#�sN�[�RҊ ��\u�ec8V�<�M�w����;c�	�TI�fDVKofR��̋��DVfR���&3~}6Z�����Q�b��7<9W�s���U���e����F3��`�&)Nc�h�SU�oyr��I(�P����%f��;�բ�܇�W5y:�0�T�,s�U?/��v�3߮�fD���-XW��?����if�R��eE����*��-���G
X�q��m���n�e��vlC/�<@1��M��'\�q�Y W�C���
��FG��|b��������Ilղ�9����Iq�j������s���[���'��m��	Q [5D ����5�JI^ʽg��j�?r�l\�>��j.*���G�C��m3#sTUl�Y��}�Q^��,�WE 0������g��6�2Ʃ�T���+�H[5-!X
��Jƥ�	7��.��w1��g�҅iS��������0�Ͷ�d���	���|�J#����Y膠 �-t��j. ��fl߄g~z�e0՚�&�a��*(x�*:u�(
(�룑����}� v��a�w	��f[[��
9����M�H���"V����&�N������Zg�xv!�e�\�i�e�gC�.W�n$�����S��:6� ���r,-�"Pl���ℿ�I(���ʤ��hd�0��f�Q)�%{F��G�']N��D��D�����]��>et������d���N���P�vWz`��e�NaYA#�gm`��Nb���Z�[.@�'>{��b=����28D������sz�h��vA�`���C�(�=�3w�?�|�_I����U�:_7Q�уQC"c���� 3���8�B0�}�ԁw@HEް��*A�+���	OHvU�=�F�jQU�='lN���z��#��{�(��1^�+�S�Ŝ)����7ȡ�]��⿗�!�lGz~C���8���3Qi��f`97D�A�I��~�1#�|��"���A������{�G�ڏK�.����_{���"�=U.S�)����L��p�Y����r��?w�Q�b�Il+����k�����F�_)W��>kD