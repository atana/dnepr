XlxV38EB    131f     4ba��b�NTC0��8�Ԭ�<C��	S����v�>��oi�ة�t���u[n�r
8����֩c�1y��T����*�8S��=!��P: �)�jy�bJI�@徱B�D�FE�o�=�f�=sexiSٗ~��׀������1�N_3�.|�s�ވp�/�&R�p	l�jOpKחm���!��f������2w�-�t�R�h
\O�rY�n'���a&XXlj��vc�D���F�1���J7jhd�ā'��9����Ud�&��]�
c��/W�'���@�	��-�G����;)�b�a����z���ݻ��N��������)��7���Ζ"ʻ�O�݇{Ì���.��m퀠Dl�%t���m\
�9�������d��j���U��n��������/&���5�GW:��-�C���~?D�WO��k&�h\:���D����n���mh����2�v�^诱���j/j�ie�5�m��EG��#=�r�~;7 �rH�Oi��C�9�kYb8�X6w/Λ\�Z���V�o��j�m4˅��E�������[}l$<8�5�(���=ב֐Q_��4�)�Qsx��3�̔O9������|��Tw��זA�~'_#ݛͤ`s��엱�V�tk��Z��{h���B�*А�����FPR�,�C惴L��B�B�d4��ߕt_1�����N����LU�tW��)��λƜ�`������S�+�t��to�qK�gq�Gm�1I|j*C�v�*�[5{��9���S�%�z Q����IT��W��&~�������^.v��7Q�KG�6�q�������Ў����9����)
d�<�ߐ�b_��O�(��`�s�5��tUW�@�33t��l6���o`I� l6p��bЇ�|�
���"''�$Y^�Rq"z��q��߁����t|	��b��7��N-�M'��ǐ!2��۫G L����r�f�fE������e=�G��")7�`��Udm(����������:�=F*%�&-�و���swP�?ޗκ˂�������N�Q6^o��/q�D�!z�#Uv�~t��Hq���ji"�glv�S_D��Pɥ������ �}jta�KO*��񲯌P/������LlP�`Ȉ[Y�6�`�2��N��2�e��JR�cgG�|�