XlxV38EB    193b     6a1U��=)�x@[	����TS^=��t��ƚ�?��5�h��Jzo�E��X��MH��5��Sm�U��w}����@��,1
���)_p����3�J�I����ՐW�R�V^?JK3��.A�����P�5ur��V�KR���L	��$)<*�c]L��é������q\����NQx�+jW�ݿR#Ɍf\KD-}/�G:@�Ьf�-ha�&�=x/."N/���<d��.��+�t>�=���J���CJA`|�33�P0�e���L���~H77&]�I~n��W�iO�R�G�p:�KI�f�|z&�CgU�b�i����2�f����HdZ7�+����_��_j��(�-�_��T�ξg�:�Ic�O�����Q:�(�q��v��3�*&h���S k�o*��!�?���:��A2*�O<��3^^��C@p	�ɺ�+EYi:������)������e��9��+
�?v20P�:��+b���;���ݼB��E0@j$�� �:-���Y�IP�����wxȽ�(_�ϩ�:jN_Q�f��9�`�i]��H_�����>3��H�+y�CI�+i�k�~Xlxs�<�g��9\`B����8m4 (sG�|{��_�D�Q�S�j�
�N�/>����s������2��xb�Mx��G����i�����$ 淃cb�mZꤦ꺃�ŃgW\cL���lȋ1�Z�c��1 A�}����nJ=�o7N�7S!�� ���4���մ�0��� ��� h7���y\Zܛ�K�<�Z`�q��)��K��2��?�K��[��V��hhk�g]AF_�� ��]^��.^{����\�V�˲F&��3��%&'|�u������E�	l��b_�P��43�[�瑁¤ �$�4��V��!y����qz��
�[W1)n�~V�d��L��f�M9�E�X]VFx,�N�l�t7�/ ��?'�a>��)��X"�C��{�{�w>����	buG-
J�t��G;084o�u��G��� #��$�zb�H��AY()B��ê��?k`P�t,���J�c{!$@�W�1���w�o��C�T�OH��h��H�(}�!U=��^X���MZR���G·aC�hӉ�"�q�5et26]��Rg0�4�
��2�7л�H�)M̊��6�So�.2�,���)y�I2`n�k���0�Eܢ�	�����׳5��e
�^0:���-�	_:O��#��w��_�.'�˴��o�^� �Z� ��GBe$L����̑w��6NpN�Q�W�]7o�$����p�Y��X�G#i�{��:^&����^%�����a�Ы�L��@�?;L��6�;� ÒP3���u�`'�vT��za&|�Ж �C�MFʳA���!
w�QAm[�t��t���� J���)��k�6��VM6�=¡o�w1��������#�1%�4Qyr�î�=vGK�r�' ��|C8�����]ݒ�&b"��M$B��7�Q _F'Jkk*����(+�H^�ǒ�����2�d�J�5v"�1F�u��2�����	
��6�Zzv/]U=���:WP���tۂ8�f7����S�M���@$	y����[[Ɂ��^a��~����]�?u�ˎ���C2v�� =>|�~p����	�"��\1�z�~�a�