XlxV38EB    3ef4     ec5��^���Ab�Kc�y�%�xx�Ԟ'�S��F����jߵ**�$,�l����|�a\n�?M��A��0�l��8w^�Pgt�b�m6v}rf�y���w����u��8P?� ���O.!cO�G��_ �\[�df/����[2�6�B�=R*�V$� ՝����'k16ɻy_Y�	���׹�5p񂏵SP�X@Dh� =~Y؊l����oin�>ߝ�O�G��S�l���kN���޵Ԯ��6'�d
�`��Ѯ�2��a5�Z�q9N�Љ���s�߸o��(�5uT0�ϑ4�|��OH�0 ��q��nl7��X�Iԇ��N�w���6��H{,�; �kC�<>�������t���C��+/KsBXu�?�#������.Mv[L�gs<�a���Ȳܢ�y�I��������?W���M΍�&aTî�s�,����������rT��CPi�+z�d�.������_�t��4W�,>���X�_1F<��p���o��w�s����e�7��l�bڒ�m��FHԋ��U ��\n\�H��x�u�/�8 �u!Z���=e==)���[��1<���ule�"��yY�冘΢�z��UB���:�-�$��y�3��m����V2�����#|��Wc�~z-:�lB`�8YT揹&�����;d:��������Q&�L�JZ�sf�F�[����~��u�/L�wD5����Ѣ���F՟	�O�1H��Ȃ�Sa4�Jr��Ԗ�H�|O�^��w0�MŃ�*��9��T�G
��g�k��.�@����7{�&Ol�}h!�,q������p�����p^����Z�����(룗֊#%��MTw�z��g�� B?c%�y�D�Űjj^�%�4L����aȹ,`�'�23Rn��=��uV�7?+/�4�}�Q�)����+�ͱԇ��� ڨ;�D��Σ�кQ��U�n��,<�1�r��<UϚ|wVcr�J�p�v�Y�'��"�%Im�q����� y�g�gf0E�[l|r�0*"ϱ�q�R�焈�N�����O��>�J��>V��O5�H�ķv��$1K,ز�6�f�q7u��ǚ��y��ݏT���^-g�kۓ�@ܒ�;�=����r�#�i�k�R��I�i<^�.��b�m�Ip-���/�x�-"E�F�]r9pM�;�3p�˖����`k7w�g��[�y�`H^�!m[���(�����>3��z�C���j��%dz�y}7��줔jf����@=�q_EGG^r����G�gF�5�L�P7�i�j|P�Npq��v7�P���,�
zDl��l�J��.�l����W�Y��q�2�p�܏K4Q�j�����d���;���1n$�M��!:	��9	�/��+��$��c �D�<��w����T�y��e`�kΞ��K�'젇��*�&��4��"���b��T��֌fo�H�k%�Lkd� �}�)e�sN�
���l�M��|������ƨ��2�o�Q���-Ki�c��ؐ��%�Bu���8JZL��I	6,y��o]��,�E�.�M�Ê�K��cXs6���㫢� �6��׹���LuW ���S�H$V�LM�oT'6��ܛо���H>��5Z.x��21d��c�8�JH��3�cU��� 2�;��xڃ5XC*4�?1�֜��t;շ�z�p�:j�<]�{I*Oe'�*"��9�d��a4��%������1`�g��|����Іmn��8��v(���>�=Oh+lFI�ۜĸz8�����T�k�e��`W���BP�:9|��ǔ��=WS~���	]�+�GX ����7s3PA�_��Ȋ�L*����&x��h_;f��F�O/��4�4۷47�#К� �F�#K��J�Z2�J%nP�!R�u'pZL�Y�n��6���	���D�Ri(ZpJ��?�#��zb��K�Gjj*��*�^Ok-^t3f��Έ�,5��H��I���-��#�Np%ʍ���'�Q���Y	R4 4��1�N�OĩGx�_�T��$��G�L���k�ʖ�"F:;tϹ!�:Q(3F�aWi��@	��@?D]O�{Q�	MI��xܸ��85����Xa��iu�\A��������H,贓
����C���?� �/�q�+�Dq�fƪz���=:���{�w�N�6�~�@�f̲B^*]�+*�q�r�8�T�M؇>�M�:Y��:V��Ɵ	�`�q�qE�M����_���'�)��24A��	���������Ы���D��z��`�4ō�Z�
+��iV3����No�z��7T��7S�?.J8��_ey4�$������w�S��J1����˅;V�KT�#P�䶽K��P�B��9Ks��0ځ���Q?��1\�u�(�]��,��'8�6��f=�Op�D�M�#!dd	�1���)zu�SF�2ӓ�� F��Je~|>��u�9��×��̟��i�`n\E|u��OK��\�9 Vʷ��p)���p��<�u�b�
����M�w�=+o;��4��y�uU��u�:&�v_n���ț��'J5��Fń2��C��B)����6WC�]�k��Y�i?ʠepVd��ż���+n�4Dg�B"�R]��F���wJzo_����a��P�Ziolr�Y�.�Z6T��Ye	P��oX^K~}�HOt�J�Y���~hŠOj� G
����!Țڰ��%Jj��[ ��x��^G�1'��u:Ѝ�tAg?�'hZa���V�u� [���H��p��E�D$zQ!J��ɏp"A�:W�ɊDb��Alq�\!{
	�L��˭���{y(��_��c�7.���GZ{0rI�Icr1Lis�lo5jg��}b���~G?8����m8��$�	��,D�Oڨ�`ݫe7� ��%������:�J�/8J߰C�,kk��&�b�Ⱥ�����P!~_U�Xc@eM����s�C��b�����eX;+_f2뿡��W�/�CŔ�� Ogw���Y�;m���N�%1['��O�ۜ���ݽ��[� ����y�����d�{�H
/�9�x��OxŸ��EF@�'7��Q� ""3�FC�qUq�:Z33{Mgd4�3דĶ�.EL�|U�c��r:ͽ���(��ڃ�:g���Q���x���I�[L�)�?�䃒sN.����_�~����FC�iES�[�d㜛���Y�#$d��=���,,#X/�O������?�:
�����4g�I�Mz�84r��`H<@�ě���m�0	�ɰl���8�Z(e1ҒB�@���i��b�F!k�����?�ȱj��1��q���e�2BM��2�E�exgM������F�����º�<sJ/�A��߽rOc�_�,�2����姕���/"��#zV��;i�!i[����:W�=�k��Yf��a�k��'>����-�)q��P9� U�o/�g��U'���8_�sbu���v�-��P7bZ���&�H��!��TG@d���&�S0R�Y�C��H I��MG��>�Ԛu�|@�a_�'.��r��ʉ��q��C�|��C��	a<1������F��Z�2aa���XD�<��v��v򢂘��=zB������䎿�-䁂��L��\��2���ў:��/)���{6A:��c��,ڴXT0��E��Z!E�Ccw��0;���O�	`�T}�h. �1!�