XlxV38EB    359c     a1f]���y�ȉO ݛ^��g�i��3K�r�އ!i`Z �ђ��)-pM�a���P��iD���j���+�db��.2Mu�c�� ���ߕ��āguu����ҁO4�)R�x ���]�αo����)�6��$[zے�7�l�vS�`MrlQ~�wO��q�5�c**��("��scr����e�x�0a^H�㛶!2�X2���cVb��w�գ�ޖ�)�/=U�2ZX�'��x��p1I<���'(њ^]Nwy�'�#נ`P2Wť��U<��z9�����{#2�����||���.�eMW�Pm�7d�H�q��)ܽQ(��fE�*�ٔ��|dl7�(������I�`�݉������svn�ǡ>wqI׆A����x����@��Ŧ��nCp��~Gy��zֳ"�ߎ�k^��o��ظK�h��y?3���a@G5�82D���)4����o�M%w?ed�S[���p�ꋱ�\w���wBNX1�]~ǈ��÷�60?���;|����?N�#�;��,�Q?�`��r'iz�^�	��}r�W����L�=�,&�%�%l�0
���R�ѷ]�V���_p�V�<}mSxPIW�R�E��r�����)9�À�=�?	�& �T8?Z�w�������yM��#�b!|�%�Y�b�y���z9=����)]2�ڳ.�[2��kUa��C{$��!݋Py��n)	��$��RhlMl�Ӻ���� ~��$�]]$���K���f !���IӚ$�����6�M�9x��eo�G5���P?�-�\l�k���X8o�`��n\��6T`�3��h���/$t�i��Q��Q�Zd�lb�F�	�{;"�F$�TjT�\���6��`������YC����˸s��3�f늉���g�Zi���-(%.ֈ�wO����;�v�6�.�����>�O�\�L�5��iN�A<PCH,���Ľ�E`�%�?-���� ,���0I!*�%0�iҥ ��"��}��Q���RԄ�(}���2�J���5���%�ӑ�M�����畴7 �VD���vcNK�<*���k���D?�"�u�hY?Vų�nY+_]����o���_�҂�M�֟����<�MAs��-�8��h�]��N�����I�q��C9U152� ���ݩ=��)�1�^M�:�W�{V�,g��n��'v�y�'����5�3OԃS����*b������?*68f��&��VU�Ɏ�"ON*B-�zz��|#G{4�PX�rr������.���)4��;����N�k���k��Ll��ϗr�������7���]��/��aHr\(f���b��}�ŀ)L��l	�r/�?Gg]^m��W����Wﴷ&4Fi����j)���I��:]I~f�n��D���!�RJ��Q�)�����"F�����D;�k���b��GMmr��N`B3�4�<��6���qIP������� �������f�C�xEjf��W�9(� 
�D@�s�':g|Ɗ���`��=���0Z�U@�����
ܑ�N>]럄z��M��!78������;�Eİ��$�@62�͗8���1���'�u��C��h8���5(��c��?�I#� \�9N���3��~.�GU��������¥Ďidg䘕�!0p~�O�L��Vc�n�F�<X��G禐���\j�ik�k�n�LX;ϊ�Y=��U��J�u����Uw�ε��`�+�kT��A�����[C��(�LO��t�X]dƀ�\E(� �E��;�46�3�]eRx7�ۡ(C���I,|)Sy*oG߀�LcD�7d��73F��]�ȳ��M�x�j���֌\$C�4�>�a��C��U���P��o��sYd�����Wj�H*/��	U��Y���[Ww��K�K�sp���>^���A�;BN�!09	���d�9|��Z���άT�*b���6ǧ�4����%��F�5���v�`5=�@7��4C�X����ESW�MG�>O�Ib�a>��-V�X�ty�W�/�b5ʏ�ӌ2�~������8ߣ-.�� �,�;��ScW8�W=c�U� }�����q1�xG P���o7���˴$���
�bԞp��H¶����5��7�9�� :U�j%�
C'�& 31MDw^}��I��f�����x1�99��	�4�b��:�c���j ��5<�HQ�ΏI���H����?��疌�VUA31���@LNU��-#|{��(��.�t���a��]*�x ���ݥ�|�.K���W�S3��@�>T�G��������w�Σk*o���ڭ$��ʖ�ý�9*9)Ѕ(�$�]�w��������aap_ �So �ϕ�-IH$�Y���H\e�Y� ~|H��5 �rf�@6�!�T�^�B	�~�������`��n ̮-lٝ���"�B{�ͪ�AezkW�(L�/�Y<0in|��/�GC����ϋ��B!��>#,�{<6�5Kx$ ��ܘ�Z-r�eP���e�=�