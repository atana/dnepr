XlxV38EB    1c64     64b�\;"F�j
4N�s1]#�V?����5ྮH�O%�Gm��ADڤ�VS2��@סaPc�S�7�0ZvNł2Z������{Aʁ������鈣����($,k��t;�TlDH[���J�{LA��y��OwN3�`
�������|��|a�$S]�vX�D��1��|}�ji����yY�5�&E�.�c�9-�E��׭�01��%i����/x[1�n�Ր\���cxQ��`�.@Fߡ���[i~��5�Q���5ˠ�
�Փ�{I��[�2����f4<췞4����5�B��g�{�'_U�Hv�2M/| �������'�B@�G�9���!�:F�]}�y_W?Ț��D4u���1%x��Okb�N"�K�g=0r��*ey�'�B�t<����ė�֜�ǑW��8(����K�$������(���.du6���;��x�Y���p�1;��@�o�(xc4�N�>j�����l P�7�G<v�2��{�O�)+��׹��:o ��В(��[s��epb����,���X-�vg����^�Τ6֝u1��������?Ʊ���U:������sBE�4�"�>�t�R�L�&����5�eQ`�RS��,��8�~��KZ�c����]�rR��L|.)t[)y������.Z�F�]0�*���g�>3����
�d>�* 7|�J����y�uH�T!^g������e<H����i���B�kX���'�R��{��-�!O�cIq��ڜI�~8��;�ԋ�9��>���pìz��1X�� ����
���-{�C[Zբ�nE�z0
����L�zOI+ �v�箣,Zy�@�.��[
�ZO����3gj���g����We����_�-��D�غ���J��-eDi-�����Sd�/��z��r�&r�%��C�Q�:J���$P~a�`BB�u��@H���$cE�vGIWȚ[C�
ָ����TI<�{� �Tq�^�!`7�|��a�ύwT)X�&r`�E̠5PB|A�"\����H���W�;[|j��� ��J"�w�SF�d`�7���!W�Or��8��3`o��QX�GkH]��x�I��#8	c I�$ښ��sy�򮫬iOI�:#�֪��l���z���ߴ�H�>��2��2�u�v�U;_�;+QZz��a%;-~��M��Y���J=µt��+��g����>o)` �-0���WPO+k��9p!Z1�)s���3�h�Ү�$����#��8G`����~��a.��0���wa%Z,�~T(2���`76kcI��l>��N���p��V�i�$%���z�(�K�'��B�]Au��h1�HXa
l+��h�1����W<ez0�E6��˕���r�q$P����-������H�倯Ы��t��A���VR(�J�T�r�r�����Hx��r�{��L�5��\�:R
�m�YQ���*��f�,��8��y�/�l��	S��M]_6Z,0m���@�dN�+w�%��n��r��d�XE=ݵj�a�9���z�"���*����