XlxV38EB    46c1     cbe@?��;�ڿ�t�ƍ�k�]Tڪ
m��J�T ��)B�Z��r��$�[�HV�V�ى���Tl��r�t!{���65W�z �7�������\ Ye�S"��,��W70$(�e|,�ړ�N��D*&�v)$.F�c���YfP|�mT(
��q�x.T�~�P�q�����U¾J���!��6�G@J���zWK/��W��a⭎���-�y#$@Y|��	����� bA�WK��K�޶y�L�������[.C|���E h����!������\8pJ=��ݐ�&n�"L��u�"��&L�TG�����ƻ
�
>7���Z����b�c��Z����3]�O*�sS�
qT=@ľgJ���F^[��L~�j��l��s��>o]���Nz0���c��D#L^����L<F���!�N�lL�T�;s0$Q�&~�,mY�J8�����9��L��,�s�|�ͤs�h�\�1뿪t��&+ȹ��kSI�j���Fd�N���K]4��H1�J�[ ���� edYVX**�<K���]�X\F�Ųu��`H<gEj�����Pb��@�>�_����XD�>�`�L��+�K�5�f������G"�BW�g���JkYt�>>�ħb'��Ė)��G��K$OŨ39���r�sg������W0�+�*�<68C�71�Q�����tRa���V��Gr1�����©�),~1f��ó�K�^b�J8�"RKf��fK���{�3ӾI�cL���#_�,��q W���[�`�Y��&�$��Y]��ID�ei#�R�U��u�i���P3wh������=9�y?�����8�a$5��XQ����1�%H�.����d8Ipg^p�����K�Q��F"�iX���It�i��B��ww��;�lS5��q�1,����� -'����-F���C�e}�Mє@}���H�{���i������yF /ӼVc
���x-�yp���>�<�d�F
��@7Ԅ��߃��֧t�-aU�RpM��;Cqj�W���h��w��6`��'"*mX��0����A�]����s3BP.d�y��L�̏��?�J�NX���!�MŤ�4'0��<�	 VE�T8F^��,c��l��M^����0J9{�d��=P�6.�#V�q���&��sƹ<�q�V���`ir��\��
Cɕj:x��Q?�LQ���m���J�=�7��{FF:߿�;YSv`[#�=�[.H��k
e�_!���G���
�t��C}"���]�]��W��[Z�D�ٺ��%����A�^f7,�[P��<������=�=У7��ZA�rKC���RE��j�1!�o_X��X���+>�5ɖ>�ڰK���Yp8Ino�u�죐FU`,aI9q������q{GN\���z����B��B���ڏ�#�L��[����应o�����������+j̜Ӑx��F���:"��٤Q�s�z�r\��,�e'}D*���1O���p��D�jj�E����K��@,X����0|���y��O�m`�	㖖q�f���p��k�Y�T7n��5�ʩH��6�R�9�$����N|K�;��m��5i@��!c����*��S�ق� g������r�3�-w�٘�����{X
��g�S�>�W��F�c���z��"!,���/���>9�?��f#w��=Rc%��I�G�YǤ�����k���a (��L�A��.q��Y�.���3��Dm_���/�=ܶ��$�יfjS�4��Ԟ���*|��R�
 �Y��LM\r'�[�0UmĮa�Z�.��L��؟�݊�x�!��2��S	���*�fn��sd���41*qσJ�:�z��z+Mi�s�	�c��:���V��f*n��u���F��Z$p�����R޳�v轟�T���HJ���|���O%s�܅{�3a�J+���I�Ϛ��ܔ�(A�W�m�xe;� �ح>%��9ź�i6S(Ly!Ɠ4�>U�+���<�
%��Q��++�=I?Ó��{�|4��&�5W����nT��V!�P��t8�5*@6�j���~����\�*����(U��M�Y7��6�4�QK5���Ig;NX�gƎ�;���LG䂷XK�^L�	*n�,bZ�"����_�a�%m����nTn�&�f��8�h^�= �c+�@��5{� ��T��@�6 ��`w�>�`�$�Ii؉��Z]�ء�V±�T�1�HRʙ���V�t���\~(`V�
]l�/C��NdZ�cXG������o�u�Y	��Q���{�y���:,E�YHb$���F_0�D0��L�?�a
cMs�8���F�6ħ:'�,`� &���85��nP����' �%���#�) 3x��[gT��[V1�Y"]��9PncM�ޚ��~B����A�XG���{�f_��b3����(,O>�3T��� #�?SxlrO��Ek#�=��n9���:
	Q=0�]�)���Ѷg��:���Ȃɞ~�/�	��2x�'ɪ�]$�8��Ci_~��<��Kԕ�m��2}Y�����[�7�XcO�47�w�G#��u��]�;��]v&|�2F�Q���4�*��W�'���ʀd��w���urR����-��
����.������(x��ÿ��oU�LdYz����3�1��J��<�Gg�.�.��X&���y��\�����tI>�dfW�-Z�R6L��/�W9"��ײ�5+����nQI�e��R�
�?�-�V/*P\[P�M��i��&��4�]��g(쓍��̔u-��m�F�u3���}c�����q�3��a�{�U]K���h�(G�ʟ��)9����ƃ=U�֭D4/��O�'،�|�[��xxh{��m�Ԧ%��85�-���7T#��dE���J�T���yD�(�:��,sI��;eggc�v��Wg�JW5#���G�g�Z����Pʆ�o+��F�Y 0�)��%C3F��~D�����c;�z��&�-��l�k�8㳜C��+��V���Xv������E��$�4/�;t=��ti4��آ�C�`#�v6��n�}�3���[�e[��U�5�Y�z�[A�;M!�EF��x��l���*�Sî���kg�}�u=P��d��R��\��1���� K�h�