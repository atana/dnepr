XlxV38EB    26c2     860&`AP�f�_�6]d�7V,�x�%?��z�k�gqx�IE�@��x��ʦb��?\�TU���H������{֒�����#��%��ֺ	�o���O>��|��ԈKKk�߮E����Z����W4��t:��[���e������h��'&�k<�*�|����$���K('*\KK~ǈ$)5�3�u	%�8���~sL�(�	}@kD1� �sN3&�E�(��ʓ���W`���28���y�gei�ӯ�|Sl�E��d�=\
Mo�|k�*���m"��,��@�-�м<�BMUy��6/�I&RX�`�ˬ�Jҵ�`�ʏݮo��o#F���Fz��A�ٔ��o��*�Ӭ�l�q��&b}��X$��9��UJ�+��Z��	tsN�ʀ��wel�-qimI��*Y(�%��nc��M:=QeE��U���.��K� ��v�V�|�-<ǍD�%)�L�����l�J�35f@��_��1\#
i/��{=vQM�YC1
BEn4��t��m���c�DTh�02ȉ�S�JL�&O�.��ݝ��'-��0R�d�s����o�<��o���z��.$v�r=�����S��΀u��H�9��&k2�����j��E�ôg�u����&��I���w�}�yi�'�R� �PI�"�jⓤv,-�*N�Z���8�P�
��,�'��@�ERG:�^0K�����,F��B̒Qw;�7#�ҏ(��eπ�Y��D���̯�ӝ"jk��\���udƎ*�C�)��;T�48�E/n /��h7pE�v�yÚ��+I�Č�y��ܧX�.ŮA?B����a�ؠj*�ڮ��t���Pt��N�4U�K�$��Q������"�����X�k:Lk��L|�/z؊��������i|���U�}Yr.�_��=燺@Lb1d<ш�,X1�l�)ՍJ)Q��m!Yߪ�G�7/-u�B��v�� �)�2l��/��"�t���K��q̟šR��*��$���S;M�8��-�	c'@��9*2.�l�w����P
��:�}�r�א*�Pw�?�O����ǧ���<A����F3#ԣ8��(�z�;�P×�]��S�ɘY�Vo[�4FJ$��ĘNC��{��CF��\��Aԅ]Ǌ�|�u�J$�LI3����đVڊ�ԤCl ����0y&�Stb/�w�IW
����o� ��4��4���b��U����E����.�G�>ѫW���5-�l�����kJ;�h�-d2����x���251��W ��/����_��S*U�;���ߩ<�5fH�|X�^_񂘆G���RO��_Y�VO��A=��)�)�
�˾�{�O�̇�E�"��U��i��Sه��� �������h������`�Q�p��GS]�qne>���zQ~��cXﱽ��Y�)"�����;16�W��kV`WPX�(ś"'~Hf	Q������ņ0U�`��6��}�d�e{�N�T���M�R�a�A���O9��Fz�U�����&
W�-�AUǽ����'�%���7��eZU���=�6���8�1�����U�� ug-�U��[{�'�
�  <�l�]��Ր����I�]k(-���'�O��:�LJ���ؖ���$Ts�ࡥ'_,�d�� �����^
�鬣w\�;�
@�UR]|�/��J��k�}�҄=b{���YAU���9�L.����z]� ��oODvƚ᪸*X�i� �+ż,�37���d�:-_��!�OT�|o`KTrr�5��ֆ�YȦ�+R@���?�m.���G���x������p?rU�ʈ@�3�e@�͋zJ4<��v�8��T�<�Ջ��+����X�y���νj�tI�3�x	�����p�o�Vڜp�@C)	�>58�D	����q��qT������Yy�5e{��8(�23�"0**<��]����_����%��[6�"�д�;A��S�$��tj�̭wc#G��Pc%�Uc��N��t���A�� =z���c�}u�j=���^b��('��
a�#�<�֋_e�z�n�h���|(