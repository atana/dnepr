XlxV38EB    13ff     4fd�)�C�y¿�]�kh���ߢ��G�\���&�*�#`1����R�q����Z+��mp8n�:`�FhWû��`|re`:� '���G�U��>4>«�<����E��Bz�<8;i���u}����H<�����{��[Ӛ�o���*a���7[���J:%t��tl�Y���RF��r/�;�g�@�1�&F��`�m�&�����n^S�B���)���`�Z<��I�K�i�����͚~6��^+f�hn�����@Yj�Z��P8X{����p�R���h�i�:�!
E���b{��L����������Nomq�����6��6�������5_����K��`�y����Ǳ���6w�$�0s���<@������` \�m�H $���ZB��7�R>�s#��[�/Luz����ǜԢƳ�Ȑs��.���l"*,]Ge;z�������%U)?AN��)`�F��Py��ð��E0��}QaUK�yD v�)�x�Yx�xP�\2`�x��y��'�p@�O�A��_b��9��\�,J����ȥ�8�>Į{hSl҃��P���ǻ��άׯ��y/����&���� ���7xB[5�����^�6W�^�;�N�Jz�t�$��E�޴���P��h��w�׺�2HV3�Q�Ji����ɼ3�@�X}�c� {D櫋����JO�A��Q� �%,�AgrU�g�~����P����&39�${�..�!��A�ުpj>K�2Ko�L��O�e�Ʊ���!�+�:Ƃ�=ˣВ�8-�c�1�lM�>�)���OCf�!sw�1m�q��G$��L�N�?�[��@�m�1�Dّ%=o�f@G���9<9Nk�[,�>�����SZ��
O\d��L��� ���v�)p�����LM���XQE���E�բE׉u ��Q�G�5�0�@����V҄�	Q��"�^=#�4������6���\Dsqe˘���Y`sϠ�zı
��-�@�w����1�Q��ƻ���x�ɀ�c���"p��k5��4�@�a�x�&Y�^l�^FPh� �ߵ�D��[�m�&O��'���s��+��6�Ы��$nb(����+��XP0a2�KD�g��\�):T�i�@5�/t���W�1zG{���!���v%Ϗ��KC��>@55�����cj>8����Q_�_)w3\��4���XZ��~�\���4�;�i#��#I��֬5�8"Y�$M�d[~n��<�T�蠘,����4�p\fo��E��	D��Te��