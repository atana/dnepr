XlxV38EB    4418     cebUН�����:�&O���ɥL�)q-y(�Ͽ.Wj6�_1п[6�����Za?�n�����`8
#��˳ ��KS�(��?�##�3^)��&{��~��k���6��Hb�u���
B�UDSQȨ���I��g/;h����:[͢����%��˪+��L�x��V�*4�Nօ����;\���-%��ZGY C�yX-.wk-���g]�,7�����Y�_����7�Q�����$�u��U��K�����jЅ|P� �F&�<��A�� �a�I�w��!�TS-��@ʆ���C�ܦ�,u�?��3��ڒ���)�tx���C?s
����/���_bٹ�^5�dp�s0/$!�/����������ť�=oXK�%�խ��N�+]�9�$��pa@��ɱZ�и��8���΍{'&i�~����it@+V�A��&�9acJB�ҫ�8+�l���"�3���iA?8�^�^?y�݂ͼ}�T k|u���HwT�I�~J;�,�o����/rc�tE�
)cg�\Q�b')�f-�5ث�D�V�ā������I��:ڞN+�.��<N��W�~F·"U�����D��;[�V�\�v/T#��}�I�u�L�:�~�����;�pC5��@6�괠$�v�j��"��ג"ud�*��δ#P��y����\�\��z��ӸEѕZ��b�}O�s�rܳe1�L����+E&f�]�����.��w�M��*!Ģ��g?dӌ�;�?�?j���U��J�f�IYQ�����#VF�Ǔ�Ć��_��
�� j�ʉ�n��Sd�Њ��r�g`\(��@� 6�!q�@y��u�k���1��+�
J����ȧƼ�j��IT3�ĭM����|dA��pˏ��3ëط�����n^���k�	��^�s�Q=��w��%�2�	L*��`p#�S�lmZ�R�/xu�	O[�O�9+�
�?1~ر�w`�hؕ뻁�fZ֧V4� ��T^>H"4���%Դq��sg�ĸI������(Z]���A�<R�[*V�d6�f'�I��������O�7	n�����.91�Wc�D�v����s����yd�C�wnɷ�c�2��K���TPz�T��]�>zߴ�n��ղ/���$+%I��O�tJ?!��Ũ�x�hY�f=�{Y�ZO�E���X�B�rg	+�#[����|'N@�.�Gn�B��G�YI��x�Cg�~qs�_�f�wMRs�ݻ��������^��gO��Ε��&���gu��@�ԙE-�;��3�C^Dߴi�Ms#+�C(���F�Q����%/�n/'�࢟�5�����w��"�&HH����i�c �5*��
A��ʹ��E�^���$Ju�q�`��I�֔�X���ir��)o��'^0���5��H�_&���O�"�v+���`���e���3J8�V�y��պC�vk��*ΣŷL�d��(���C�#���*�j61�M��SI�lkw��ѐ_/��z���T�c��^���IΆ{$�>&�-�#�%�Y�;E'�`�ɫ� �;)o���y�Q��yAاN�O����ٚقZY�ޫ}P����N�[r�R����^�[��.w��<<1�SIb�\�BX�Y8]����~���o�X��<L~^7d��O��3����Y� vQ��$�Ե|��,o
������J�}�NLx�;L���a�/��*�/W^"ŢC�It�-EO��HA�_�潏b}I�����G�A�g��QqO�i�Ͼ��
�ɝ��]iTZ�-��\C�.����Zk��[s�u^/+����m�/;��Q}�X�.l���h�l���K p�v�s�Z�b�)br}�A�cԚ�E�/:�=��:��r��b�W�g�����|� A��s�	�&d��"3������Gc ���vdpfE��`��ݾ�)*Tl�ۭ��zxn*զ�.n��ϓC���=[�a��������{p�9�F�Qz���Z��>༓�u�yg:E����d��^��R�=���Vd��n���ͭG�Bp��ƿ ��{L��E�ۀ��Z���S
!�`�9+�H:�]��o��R�A��4=���{���UPG��')�����A�y8/�}�%ϡ���7�󮬥E�ZJ����N�#X�R�i�p�/#��8�]>�S���fD~ő�tyJ�wn�Q��PC3�0��h��2���r��뮵S9a��|7C������İ����M��E�l���l=�?�֒��W@��'�q��hyZ�j��LY5�q�8AQ��Ȅ�	��(�m4Ń����L"4���U�����ͤ���E���	�3�wq�� S�N��Fpm�	�˧����Σ>�� �-�b�fܮ���=Fa�_�©NwX�GI��Ƹ(�_ʺ1��1=��{*�.�%kp�}�L���h�� -���"J$�9�ox5;Dw��V���`2
�H 1^�5��OL������H�M��b����1�ʑ�քu;-�OŒƅ ����*��Oȡ�`|��H��@���i�hr�!Ӧ#I��i�A�L�D��"m�Y	F�K����(�Oi�\K(
\!@��'��vI	���Z��ra%wgjQ�b�,���i��Y�(TT����%��艣Ĕ�"����"�v��T{�\Q+ft�c7ω�|n�����e�TѿD2z�}2/@���Tp�M��H����	�;�lWLT��7)x	P E�#I���1G��%b
MX�:J7B����Y������z�_z��GW�6"�F���{8S�wi��RM���RG�$?�>�]QP��/��ßhY9*�/���x��p�C��'bR��ix�z���%"S�*u��q�*v��b!~������c�����csa��V�.��+�"8mN���C8��9�yd8�K�_2�����[�=���󤜬���TW�A ڸs���Ϗ�J߁��EW������y��CJ���`�X�&縄 ��mP����L/�	�G����V�q\&��9��/�F*��(.���}㤡��h�Q�4D`$BxF�?��d�=�:R+�МuhZn�?T��0�kbt�����t���)O�`Vr�!ˑ��M�Q���Ճ;����+wQ�����t��-ʇ���A���d��K4+�ܩ�F��a2���(iEm�_qA���t��;�y�.� g��!<uEi���!PЇ�S�k*���u���9g�t��[ec��o��s��0v�\6Q���"\�����