XlxV38EB    1171     48a�E ��6GX�"/�|ag̳8�hI|�H�(�Ό�b"��WR����Fj�?]
4�)�hjK �k�e°�'�`���/���/n��%�.���$5�]%���&��!��:ڰ���稞}���� 7��τ@�}�7��8�,*[�kᯡ��C����)�
�H��,!����;�T�,�e�$�Lf�7"�}�4k|�x�����wG�r��B�q#>�%%�{5�a�w6C`�ѷ��,�6G�ؓۮ5n�]&(�SŅ'i���I�`�N��Z^�d:fefH�@y��t���w[�Zc�.��W��05�I�/��ނm�M�7l��S�� ��̾�0�D�@?+���/����2�Aݔ�|���p7}�C����Ց�*} ��e�m��i,�eL�8V�!6�
�Kh�6�wSy{Zg��,⎵-�-!S��vqc�4#y=�U�u�v�#�7�v=(D=��R��F�9l@���F��$~\���N����`�$��>�B�_EKfpB��#M��Y��P_���V&ωkZ-űa��][����-.DX��J,Á"�4vƧ`[�ⷜ���;o���2� �u-5���~��Vh�?��E����b�*X'qi����&�8��	�k?�sm?ʮ�%7.LnW�\͌1�~3\����pѮ��A4����n��7etF�e��&���"��i��N�6r.�N�����_��q�H�hʓ������(�g�0�Zmr2�S��Z%�u�h^ۼ��;1P5��X�,W�7�T��N���Py���ўI�;"�v<ØVo/�	}k��sX#I���o����W�s�qDŔ�.���r#���1�6����@�MS%�����V�D$�?�J�@�u?|aH�%ݫ�(�V$����*`Q��M�T5�ɛ��uF� f��v�Nl��"e	��#4��.��ʮDH���=�S���Ϣ
4ᵕEFXe��s=���;����|c��afA��ޥ�c��\�Hj��Sd�xr�ā�#v��yC�ˤ$)[k��U��3��8�~S-=��C�y��b��esŤnHb �^OI�9ā� ��ӗ� 7�;B�{%�<���ʈ�6zm:���x:��#��v������y{-غ��m�s����P-�v�`,�\]�$�