XlxV38EB    1c78     640�8��!�� ��xW�*����b���*�����ǥ�6�'J�4%B�+l	��F� "1�d+aS�
�{����8�(��Ժ  ��KiO�T_͖�X�C�L'��n�&`e�QYT�p�1*����P|	����|�
��L=�2����`��^�|��n�G�pM��Py;��䍕-��H��#i&'�>x /��{�
77�/V\$U'�0$��L4y!�e��Wk��<u�g��uD&xW֬0Q��nJ��W�&X���b�!TsH��m�^Q����O�K�h�ez��a��:<����;x�LAO7�Q����[�i_^ӏ��*�pAJmq���Y�c���Iy�%I����LJ
��ѽS�<�U�r�sk'`쫥��,a�VDj�=�K28}Z|-ߠ�9Iv�@��`O��0}:�m�g�٩aЪ���n�_^�c42��yUZ��LY}�<���i���Q�H6��HP�:��O��t�3�uR�%�����GQc����٢��vo���!ޏ2�����"��6���&ԶX�!�̜+ʒh�~\NHv�Q� `�h,�_C�J�aoZ�H݁т`5�L��j��02�Cj������S�k�� �ʺ�T�(v�.�����v��ҥe���!L�����(��v�R4�O!�!���d���V'[�&�ED�'���ʣ���,�q�'�����Zm'7 ��7`F��:��+ad�K�7\%��v_���/'B� ��������۩���\j3��	/ؖ��,&1J��wd�;��%�M.����R�c�F�WrEԃ��KG,R�|���m5ar�m�EJ�ֳe�����k�Ez�!���ͪ��k��`ƺoM�P]Y~"](�a�RH$Z�5�ZPprQ�0�P��Xw6�	����8䰟���?���&��G�����`�	����#�<����6���'�6i�6���Q����v6�1W;z��5
�g̴��Լ�1��d3_7f�~)�7N�vuG�/�����������n�w�e����*�4��H��JW��% 0N��~/�\fA!�BD9�2f$�0��a��OM��sh=���5P�p�^[�gc%��?�v{�]�M%��F_B�<�v֩4�]5{ty�ލ� �t��I1cb��եY��1��<���.�E-����b_ֆE~Y�O���\Z�����m��21���cq�T��Ͷ	��R��';w��>R�
O�����}�ia�N�"<�g�ˌc�#R�T<�;����7�^��.HJ�f�(s\����i�3'���x��@jk�)綛���]E/j��@DA���ТG�C�\�n�ֶ��#�K��H�TO�8e$��<�p�:kbyu7G$Fw/J�����VW1_�P9V�EF_L��#Y������(��i�@���;U���J� k \|�,�b����Y�6~J��WLl�5��Tk��dc�_D�L&X��g���� څW�"݁(9R���Nn�3+����HnUh>ӈ>X��kw�:�YL�2���д��)�d׫¤kj+:�u��`KF�
��5W:*�be�P&/�T`��O�%�1���