XlxV38EB    1c59     643+�b���0�	�}��2;C(��4a��
�0���_����ȅ���QW(9i����}������cW����a�c^�9�;�����d���C�6g��▐���G��~뷘݄�G��E�ܘ`�}�Jjh�N��t�Ǐ�@��c�t�U�����&��Q�!Krx0m�7��u��w&�os��P!�m�����v�>�b�H[T��+@?@,���xz!&Fv�j���3d���]�.��g�E������M�������
���ɀa'��C�f�����T�`i\(wbk�.�.aˑ&Ϙ��x�ǝ����Y��	�u�E��ۯ%7	�XP��Y0NG3 ͦ�`k�$��k�� �a1����W«:O�K�.�n���Lo����$��&�ς�y����[�9��<�]�H�,�0=�x9~�?i��;jq�\nP1�ʬ�i^�!A/�
>EQ{^�H��7d�(M�iL�؝ֵ!������ �o�_E�{>�10�n���3�L\�)��p��)0s���f�,[cx&~a_w<!*R��� �ME�����6� K)^�	$��&�k���������N�0o[��G��C(��E�a�]���r��Z�o<2�}�a? ǫ�P(�Q�S66-o�tq���0�N��
fZ�wo�ޓ���>�+�T��Ś X{��k�	�R�v���W��X/�v1�Z�%�>�Cnr�cH�l��W����r��*o����`c����H�i�n��.������c�uDm
 �텣+�ۯ�Q ��z�6�P���&�;l�)�V�&��|��8�K)^�S�y�*џB����?�"�Ud�]�z���>��>	ւ�P�0.�V�̚or��g2q��"�feuk#;����c��Wf�����t�ԁ6r�s���R���gC��X�_߱�k��{����P]����`#6�i��B�fV�$��������΅�TTh��h��ǟ'�n��~,�?���ݱn�Z�8D�w��ӷ�.o���j��,��ӧ�{ `Yϐ"uҖ�hl�B|�����o{��Ub��^�+�a%�07C���U,4k,^���l��(B�YZj�-��1)k��泻'#��0�i���`�gmK^�DB�}��3"Zc���N���a���@�+\q���{ �ㇼe*��p���O�����B.k&5Čot��Y2�6xma/B��FB<j�gT���<�P��e��br���ʷ,ղx7����/��ҌN�'�Ų4�*�>�XD&S�aSN��z}-^��cBZ�r�Ί�27c�#�X4�J�ͯx��ώ6�Ehz����w��)��yA��&Y �D�'?��_!���(�̼�ǝ�#N����q�3�P�[1b�?��u��χ�C4�K�����J����*eC�Y�hnۜ����5l��r�z�Ka�@�-�0Ճ�I��q<�,�]��>oGF~�W�r��.��̒'MnJ'l� 4�Q8n�Ȉ�X�|��+���F����y�Z���f�$����R�~��k�C��R5�&.�
`h��;w��7���ݮ���