XlxV38EB    429b     adbE�Cu�B��X-��X�����2��*�󔩏�F%��i�b�K����Uik��d���qu�L↳�����/�p��|�cE�W�Z*��L��#�Ћj�l:LN��63��x�߽oo9�Ѝ+�`�oD3gG�N�Ϲ�p�fr-�h�,����W����5� IV���?����0g��|�AXF3OoWbՑQ_]�=��-�Sȴ~-��=)ؑ�M}2*����`U�C�.�B�F��	�a��O��|d�~Y�����݁�wY�րK
��e�]\#�@����ZG�J�Q���>���/�4��2Ab�	G4c�Z\~O�6(U;�"��/�����:�;V�*G���Ø_����O��ǞWn��uۅ�Hi٠ϣړ�ϦS��6�Kdm ����\E1H�Es�Po��ђ�S���,`�02��
�st)^�!�[T�ٕB���v�iR/5@�P�����5پ�<n降��[T�EK�*>^<�M�>����־4BH��+rt3�����S��bĦ���������1��Gx�pLK=)�X�Md�G��az�h��_�wz�	��^�{�Jɵ�~U��B�]p6�Zf��%J��x��!{�"�����B����V�?��vBH��w6�~�3(�.�K!Ǩ����5��E�]��[� �A"�ҸJ9��q*�T4^���Eu����=��0���W��u��YEb��7�T`A�B�}8�Y!��sQ��/�Z�#���َr .��-)�@��S
|��!-���E�ܚl�	Uo$�� L'�(1�]��&o8Q���c�X|�`��a��o����L������1�,�Ḅ�WZ��D��~!�9K��&y� �<R�A�p:�G-6~�F���r�;���ԽQf�(,�T���avI!���ڟ�cn��KDu��^:���Y_�^|��(��#��x0�]/<[��@�<����
b+�p^Q�z�xu�)����r����$"��Z�g��Hl������^���&P	��z��������S�������c�f�X��tq����E�y.-��j��: �dK>�  ���p�Q�_�ݴ7�9�U�"%�2���F�ę:��r.���M"~�qA�c�aR� ;���נ�z�x�NȋmD3U�1M���A�3��y�A�ተKkyV����4	5�U w�ť�|�V�]���8����X�êŕ�{�͝��� fi[O^���Ċ��p2���G��eՄ���[�i��ۦl�u\a���r�mD�ᧆ*�]��������|��dG6U!�0��S���ƶ��ۭ��f�V��xJC����O�7��"�lSW�����{�5��iV�_M�N��y*���?V�w9��c�u���_�%ـe����Tv��6���#sǊ�s02��#mm� �
V"ˣ����uGq��f�͕�qlûۏ9��^��y�R�Ʒ��嗞���+��C�S  E��L�U�u�ҝ�9,e�7]eM ��.�M6���*��V�#�l�.bf��+b~ޞr��E�0 ��l�Ǩ�Z�@����Av�r.�ΨT��(���~G����󒿾��6�������qP�MZ��#�ߌ��.�u����a�[ ݊zs��8�\V�L�A����tp|�pCQ!��K�qݕ�F�e��ٲ4��b�}�'�N$ʬK�ts]������A`����.��k�C۾���:���'��m���༏up��f�u6X��t��'�`y7�s��?:��fdhEo`z��x�5t�Q�+�O���^�5�{�@Mn����O*��#��Ul- �3��`.�\Qq��*�D���骱���c�	Tjاf|�C�Gi;�Ҙ�є�J|���f�!Z����۾b����r7��=��J�3*!�q�3�#!j0mU	%��^�J@�*��RЀ�tʃc�`p����������b�uא��S�6�4;	���!�����J]K�@�PQG�Oj���'��|�r���TֱF���m���TRTz�����[lӆ��Ǽ�����*	����$b�B?�kcx����h5M6W�G��Y6����&iG=�����e�e����3�����\�*�d"�VXs!#̬$e��Lf*鰾wsˉ���"Б��3�V���-M���MV,��r�>�_�ȁ�>T�y��=��PKh�K��x)�ҁ���2u�j3� !���ѱ�����=k�o�Rbo����{�U�������>?�ڈ9�s"FXMTC���J��i؉h��о�H�^��M��;!*��1�!D��yZ�
�_�������
�[	���w���	*y��}n���s��vP%/sZd�ߦ_��W����V ��j�7�-Y3`��/s���<{�I���Cih��y�@/�gJ��'�C�"�@�a$�ιc�CSX.~�?Ԡ�O3��Y뮆��&���ª�e���Y�%�E30���G6W#��-܆�� ����mpAϾ��쿿g���a&�$����fN��#s=@ǽ7�C�|�1��
��W�:��Ŭ^2x�#�����jM���K]\9��/�}��]~����T�.8���"�A9΂��ŻThm��p���闵�9��W%٦��r&}UE#n`�m˸��Dq�Xy���彔hUs<�/�ؠ�?wXl�� ��(����$4l������.�Dj�=:��