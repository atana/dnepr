XlxV38EB    294e     962����跞��o#�m�T��[3
�Zկ*�ޕ��X]XΡ�r�j��Y���*\Ё���S�=H�X	�P�[�TT��κ����W�s�d��,�ܿ�lr�E�=���KzC�Q����t��Ȗ\��b�3�?��G�M}B'�G��f��[��8�؋�l2X��j�8IU�R<�8��	��ƴҐJ��4�-�B��x�e.�fF�Rn�_8	��|b�G�=,`��F/6IV�4��Gꄢ��2n�^�F���ҩŎ���~���m�e�UX�=�l܆Y˷&L�x���t�|)	{�A�n"�}�Bè��v��v����]�\/p|چ�P*��%���u��2U���)��GG2��Fs���o��7#�nRF�ޮ��&��0��t�MEY��4�4v\�uK��H# )���5 �ju5A��9�h�M��i7~��*�/���|j�_���)��E&�׃Q(綹�}Tt&�e[�X�iukQ��)��ں�<D9����Um�����i!%ɳ�@�o$'B��8g	�b��4�?T��$�-�tZ�#��!n��d{�_���
�K�A��ٕ��S�*:����M��JtC���ْ	�,X\���ֹ
��!ۦq�k�[�v��:��1m:ä�Yj�����?���0D�6H�D(ʭ0���!�ܹc�k�F;5E]嗖�V��Ia$F#��������a[�*2:^ba�����UN�0$4�V����ɕ���5/��!�<>ѻ�����q	����1b=��=�@�l`R�  �.wa�LY;EU��nFmn����E�`Ls��O�O���83��b��X�W�:����K�۬T�-Ј�k,K�ߊN++��ݨ��z�폝m,;��| �7?(a�1�� ������ӶI��� �'��%qbE��ڤɨ�g�7q��3��k�,^���ߢ�~�b[-%���B# �-�f^j�Xت�kʴX&��,d�'��~)����[�61���-_E��m.�}7^p��(��O.)�rl��L����~��{Iqn�����]"��N<#+�m��Pn��®T&����	���S�5�U��@J��GQ3n���kV�>�Ac��{�>Q�HoՋ\o~��?��3wp}��jh g�;�3�O��놺���[!Tp89�h7��K���9�R��,@��ZV�(+��7�oL�VdŔ�3;�L&zh��U���!�o�F��T;�^L�te��Is��D�/Ւ�ݣ��gsL�>	2xƎ��H^��oS[�q�Q�O��}�RM X�>���
F�$ce �"���dR�$�|�8Y��%o
�8�A�0�5z�_>�wF�����5�8s=D�w�sOd�
�LgY�ig��"l��p��[��1��A�XSm�e����VoݚJ��iKs0�"Sb�ߤ��9�S���;�\�>GԆ�տ�o���m�9Ү�w��M��]���7��_�"F�;}b/�Y����{1�A��������Q�>ܦ�Mp�k�f{�l�"; s���I����x9��`L��%i֡3��PrvS*��4�yPx�e�*��*��E (�F�:W��l+����\�|E8�5ؿK��'r��LX�������,Ɯ�~�$wK�!��t��h���^u���kR��3�G����?t󷞌��LwI�żNcS���E��;k�MW޻>��ґ�ZK?i<Dp\Tw���A�����o�*�S7D��}���>���|��7���\����=͠��w$g�W��h}��le�ӵF�]JP�_�ɴ�L�:��2��#�!
?([YBH*R��§���d��� ؒ�1��ֈ�!�)Z���vgi�fy���级*Tv��E�<�!�:p�H�����LɌ�)Ky,f����2._�S�F0���[��
�^%���&����� '�°��e*�!J��b����X;F�,�o��I��2��{K��"p��;w��?��_mL@4�+�@sQ�W�b�+�O�tH���F�#���X}�k>焾����P�h�9�>���]�L�`���L.�qE܇�E�6�lhNἦ�_
��I�7�l��M�5'��.�m`���U���2�Gk�3H�m�}{�ؾ�U����ІUK��4nk�L.�o|����?g��0��μ)��W���?_�h`G~�K��c�
1>�_.j֖���H��^�4>sD�U�7s��y��-yw�u��ӈTy�x�Ԝ@�S��^��.���ͮBH�]hMQ׵�e����=iI���)V��B��͡�uVX���ڇ>91���� Ya�7B�����D+��B-fq��'�T~��=�ų�{I��V�Y�ŵ5N�