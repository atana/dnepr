XlxV38EB    fa00    1bdf*t7o}��v{>
6� m�e�W�QZ��B������,RXY0yvhS�~n]�"����#}i��J4)�3z�į��G�V��t��0�f^(��(\����GH���*�
ȥ�x	�,����9���X'RF�V�.��fD�v��4��-�{o�+wi`)r�Agg$��
w���`I�-2���[n ��i^9D��E�G�j�,2D����o�P��6����o�x19]��8���JNa�*��⤘DR��JW�J��(����j��.�`��D������'�E������p���*��e}gA^�x�E}�H�>@Zr,�!s(��:D�T� ~<9cǶ�������wl. �\���>��-�٬�DݳH��C�d���b�K,n�=T
�Zq�N�A��$�z�m��.�ꇷ��,ز��7�<K�z������W�����q3�,�R�㭰�el�
	����	��f��-h�����l#��Y6hha�c��N��@t�NxP�o�s��e Bl���L'�c��RWH%�I�Ps62����G�rvK�l�/n�V(��c��2t���L%p��Wd��B�
�VM�9� `]U�nm��h:_����=_�
��~SoPOܘ�%g�{��`M�R���-貦�-o����}���{�H%Hh�ݝ�p�]��:���t���>��Q�MF��U�x�S��Z'��*w��1CXV��l��61�g\��~�"N�h�����0�OX�����T3zEkd��q@Y�G1�A��wSy��ĔP2�d���w66�m�~k �%�˔��:���+ �?��vO�_Ng'ԗ����	(NJ 	�z���Ҥ����&��BLF��դU�UF��dv�ĒqA2w�A��<�ۀ*�
��>S�#��ً�/���4����0BͩY�%��x��nOd�hH��W�X��_�7� ĵvC�R��=z'W�3oʐJy��v�-���?G��_ڶ���bQ��]q��R�C!�J�r����z�!��V�7z�oI�ch	@g�&3�c�)���F�T[.�H��'��G8�W�"�臀����Zߚ7��A7�jvn��w��6�����yx��A(P���y;�TJV�OI�B�X ����B��e�Zi�أs���x���G񉞡�R6�bc5_td A �^T�$�����d�s �Lm���6�:r��v4 �3�s��&���E��մ����d[O`Ea�.��(#s������&3"�F��*�(����&-�06o�/x��bܧ�	�o�������j9ۨ����y����[!5�
n4[IByh�X��S�K;����Gօ�R�NbL��Qm���a�Z�$)hBD�r����/�#]ח�~��dEm�?􉆢S�l�T�SwC%N�}����Fk�q��y>�rrڣTyp$>�e�!$T+�k�����4U���8��)f��N�"�u��e:��Cu_ Dx�q]��"�q2���|���Aa"N�H�fa�����"PUG����X=�l����\��)�x<��P�O;�F�:h��^;�J"�B����Y���d'N�\�q�o�I�{���=���3��'z�r��ƭ�V_4��?��dt��}��ʣ��gHէڷJf0I�;D},��q.��ls�	{|�yP��0�h�J���ۚ�u?�	 M�c��g�%t��k(`�+@��˚V���9�h��[�Ļ*��C��*�����Y�����iO/�4F`J�� G�ֽmC�&̒��<����3Z��٢7�\�43�9N(8I)FvCC��	TD~ۧ�܉�J*;�~���ҩ���w���g�e�M����@��8�V����<��ae�w�ߧ-�YR�
MVC��b���sV.i�T�ZO@�=%�l�#��g�7��}~���d�2�ĕ��$$i[�"�����|�+l*�k]k������t�C d�;?įp��,�ё%ѝd�Z��p�b�O��h>y{|�+�G/�,ou��_T,��\)��%3��z�%-MWi���O�U62[|��9p����]�QEJ4��̍v{�IȻ�KI�A�Hl��@��l�aU���i?��w�G��X׀MI�L��(�g ��*���������̼s�B��)y�F�`�5���m��slH�I��6�o�ÿ����Iv�I��b��L�82PP8tX�q#�)�Ӹg�Ƌ���9�+����H�q�@��'׵�?��/@�-C�*nM����"WksG�"O��x�G����}.����e�d0�ݔ���H�����J^OD�����_]i��N䜥�ﶕ~4��;:֋�iۏ�(1@�y�Y����Y�Vl���|�����E��WN=cmq�r�͟�0���v*pa]qPi�b����^pg%[W'�Y��yf"}3��
۝�n|��n��g��"��#���t�&�H ���E�A�+�`��]r�q��Q�:�h�&�N�h��~�GU������ct����V��e\>�J6���L��]١X*���u�þz`�8GE�Jl���##ծF��3�j���9dڋk���U^��[W��O,r/�{J���"Y����)nӧ��4�y(Ik�ёB�:�}M3e��4�A���ux���U���!�[t�![T���OU�A6�B�����r�7�_Pe4w�%[!凁y;�;�3oF�5�9K�՚(�k]����[�04��	ϱ��S�a�w���Bx�]-��\���{�B@N��*�]�����Ry!.&}�>�\V��Ϭ��M���C2��Q��&��6G�� ˷;�h*��i�x_�_~�܁,�5�QĹ���f�K.߇��o�p��DG��3[d7���u����;t���Gi�7�"��^�P��6
�R�3'7�g�� �.�͵#]]\��t �39����A������v_b��:��[��"y�:�GM��uJ��b���œ�Ρ��J�e�w�Ig/K�xZ���C*e�������O�&2tDa(�9�t�Pog�����{Y<Ǎ�N�)rc/�D�QC�Ԣ+��/�r�/MN�7��-�l� U�,t�\ ]��#���Itp�X�:v�� �C�dȦ{�Z-���aP�Wy]�\��	�6$���a}��l�v��=�yW°�Y^�I�O�	Xp���� 1������E۟��ge�U�P��Ͻ	+���ѱp�@	P2�L�θ��U2����ԛ	S7�����]�VtϗqiወD�iVQT�61U ����ƾ�;NJ�;@j���E�ԖVKj6q�QM����H0�W��dCp�@���(���{�;�!S�4��'�i
~P*0~n�QT�>�p�X^8��N܂��;"m��E�)9��GN��GN�* :1�/z�����ߙ��t�mF�g��Ee߶Н.F��J���n%�.�/ 7����"+I�p,2����;�<h(6���u:y��E��!>Q���*XQŗ�*ʶA��+[Ո�I��4�H��14GFg�GHg#�!8H��"��8��3އo�xi�n�5��iF��o ��π�c̣���i����yU*d���n���',��d��(�28AK����1��"�ޘꯝ%����_�� �q#��-*�\����,���EP��~�B`�y�>ɬ�[���$]uAF���z�%��� ?����r͘�� ����	�m�̙�l�>@#`j�oo]�䣩�9������.�O��@d���|�T�@g����I�vV-�,��	)��XN�\.�1A��c(��t�@�=g���΀:�����SQ��?�塔��*��IF��>"u '����ԵZ���_`��XS�Y�m�5��skw��ff��F��;I�-P���v���A��-�)�%�kv��^b���5��ly�5�?p3W��ǖ�x�B�IQ,#���*B�f���y���]{6(8����3;@%CD=�A]F�,�P*�43��_S�p�.ݷ�L��5�B'E�\]����5_��ƼX�y�;��$���_�)p4/�y��"Z�\��A�����Ǥǻ�|j�y02��<L���°9�a�uݳ&5�ܮ��(�i� 7�q7�l�IL�Ɉ�5��E9Ɵ>��sa��[���/yl]��G��N�c)B"�4��4LtӚlQq$P���{���I4�ɹ�o�+jT�/YY�ibx�g�8���p���A(�Vkv����z�ٿC6F������p볓N�0|����t����Ig]���o�Y�p��K�����N�)x�V���k�Y�9,�6��ܕ���/���*S�6�'e�N��M��un����"�|k*�c�L��7�e/�g����ޖ�%hI����,�J@�z��s6�צW����{���ăT������Iʇ��/���r��d�q�� ׉=��e-E�O����iqh��D��()���������(`����Ѹ�,{|���z@��4�1��j��o�.��Bj��}EC��	V�ic�=�P�0R������t=�� |�{:��>sY�xZ/3ߕ�G�&@�t�?��u	:�!�|��ʉn� }[���~>�Z������=����?��a����u$�^��'�S���LH��N�)L������7���R&W�-`i�GwvQ�m��r)��*^n���.���z&���b�����}q��0��ߌi�d��h��^�i�v?3�����/&��� �Jt�b��v�<O�|Lr�^�dj�*�l���ŇS�Z�bN����b�G�%+��\s�����j&m�����JT���~[�њEw��c���+�.��< Ғ�"��`���{l�ث����a�E�2e�"�a�TК��m�lγ"a�
{a ,|� ҕD�ÅP����T�(ny��md��B�����?W� �_�����kQy!�V��ɲ���#�}��',��)��F�"�#o�&a]4�*�3�AğX�H��ͧ�����c��:�$�TD@<V$e�����f-ĭ=�<e+˧4MƍoĻ�W]�=��LuK_T�x�;���9�3s�V)�e�܃��/Z��:�S.�"�k��<܊�}2N�L�\����Fcރ�bm �2�L��I5P�dyl|��J��n�U%|�P�߯^ᱠ>�I��ɡ�<�.���B-��7{��+��K��:��-K�6Y�]G����2O�W�]W?� �	Ϡ:�:��o �6N��@�����b
3�Ԧ{>���K�L�d�!����w@�~tey7L��XA�F��<Y�1��"���϶�p�]���
�J�V;��3] ���Do.�6��C闦��7ρ����YV��j�YH���ǝu::�k��jEC~��<
&�Tq��;�u"�x-��g,�����
�`��@n���>��l�Ƹv��y�`�T���It��
�;<gr�%����~כ ��=:E%��|�͑�4�7|��X�C�C\Z������.}y�:呉2j׺���h����;�V�dp$���$�،�?p�|iv1Q1������G`�6��\v�{/�:��͑|��e�1U_�#p���	�>�Z�jƟ#ލv��'�9n����y�_V��|*,��<�)p�Y�M�`?a.�P{���Z��at��g������tl����/r���,R�Oǉ��v�r%ƕ�����%eIN�v��=G2�;��I��`���w�=-���d�_��,�#��ӄ�H�ɹ���#2&��WU���u|�'����+� x�t���u�~�=�~�S��$��hv���)���Z����43*,�]w����� a���L�:쫁A�>�� ~����H��[�,�1�`}:\�l�y��'@�=�(x��>�#�I�@���Ð�q�#�����]���i��W�dx����*�8S�qѿu L�&;����~?[T��#���w�~�㬺�؞�_�P/�����N�v�x��넝V��]�jOY٧V^�Q�}D�%�\  �`��+̏�g��ڄW�Yw�!|aܮ��!/A�9����;�$�*aXL�U����@7�s��X�3T���ވn�1BX���KI�i6��g_��-�	�贍�l)r�q*�mW�pP��E]�>�P�� �דP��^�aiQ��]}��IF=,���aw��,V��/"ێ�U2[���-}�)$B�Aɲkڞ�7�`�Y6�tZ�mյ�^�"������+���{��ɕ=�4H�y<L�g�W�BQ�����R�ʡL��!�V��UPi�G2{����_�cO�v��?|s�GH,�`1���7���υX��#CB�z�a[9�v3�����J�j7����vΩF��+4��H��_���8k2Pz��_�$H��v�Qs���0�w���3$zz	u�̷�h\5����|��!�k��Y����7��nV�gC�[�B�F�	iW��0�=�4����<��GEh:�~��vp'�V�1?H)�X�"�l�����q���˗��c�(�����R;t�C�#��$L�<�s��9f��~�{DVP�7+��b��N[U#Kӗ�Q���m��4p��4���]� 	q%�3��d&p������qy*�ћz��	�����n���St ���
d?�SFi��!��R;#�����G��Bp[J��1.&- ˄�,�w܃.�<�NF��������-\����iF��-�9N�i�+�T�@��[ݦ{[LC~�ȶ֬x�lÒMI�����l:�E\����\;�Q�yˑQ[�	M,���{>��X�-��b>\����*o�6i+��0<_�!O/BY�9�
�"W�[���M[��n��R/!HN��㲷�J���?���%�]٦wy҈�Y�D�[T�����ڌ��nt\xI�K��7�f!Z]��DE�	��8�Gz�G�uޏg�x�w�墊�r��\�����F��yu��ɩ�9&j.	�f�@/��o_�яl�GW��ݐ}�Օ\>_v`���V0�������RXlxV38EB    b5b8    1d92;N��*�����oz�a�$�qn�@�f<�aJ�\�� �8�ڪ��YXY_�%���Pz���Ĩ}[4DL�F�t�C�鸙T�
(	�e��8�W!%)�����H�>���o�����[h�#NH��#;���趩�l�u Ŕ���Z�Q�Ԡq�� �T43�E�<K!�AfnP�7�R)�<So☨9@��s���IB�1~���r�p3�&.���}�wSz�C��,�g��T,qbu6�L��$� k�-����Y��Q����:�ob��nY|*�q�\v ��"N�-%(�2���5�)Q5ڵ�+���!�"�'zWsh� ��O����	*���G.L�i#s��3�M��)�+����*Ao�����=�	4����J"��ܨ]��h���0j��c}�ڒ��rw#7dԈ�?i�!ݻ�K���V�z
����>�^���U�U���/Y�
��ǘ4��n�n�L��՛���IA�Dy0J����DLV⺳g�۞���&�v�l:V��d���^n��ݷ�58��RL��N��N�Zd�Ἓ��`���`�#�3�b� �(�'��j��%e�R��	����	g(Ơ���Aޓ]���������4
�E�Wb7�+\�|��C���va/���ߘ�{�
��bs.�8�c�?�Lgsvj���&�q@ùPNV=N6r-�3�l|-~���Ю4���"��G����LH�B"�Ƶ�n�8�t\��1���"9�_3���6�L��z냇��/D���4�5�h��u��X��d�m��d�fPQpiLW��n�Z"&��4����mdH�H3qk*_ty��;��2g��%XwR��L����l�X�Қ�b�##�������l�kw��z����W�'rj���2�6P��p�-�e\tE�f�Ui��
<G�Fi�UK�@+�
tH�i����rwzw�K�#m|. ����x�s�bV ��ko�&E��Zv�K�����`+"�J�Rn�#�vN:M��B���i�ד[1o��0�\��� k�|���Ԅ������+�-m��6~!��<�Q(_��1;P4s9���(K�������g�q�=��ɲB�b�Ze�љ�W��������F����O~&,D�����_ּ�o�1U������'�PQ��ʇ��>�*��@��ȉ����<ѻ���M��~#���z��H ��#�.���Z��25�ºN�#EW��,D>d�ʴ=��G�W��*'w_�������TS�����֍�h���@;Π��i�]8�P��+�;���!e>I87�~�4���a[π�Y=��>²��ZD$�!-�(�d�ʐ�)v)°�΄��R�}ޙ�R��<��lY����	�a�bP���V�����J-��I�Ţ.��]�Xxc-����O�R�%pHՏP�[+�f�3w�̘�m��T�\��~�.=�4�ɚ�@�QI 
��:Ϩ��󙁠5X\ಒ����2A�`��s�k+�
��WY����KU�]�v�PK>Q� �j�|<H����#m�~��$-A��	7�ph^~L���䁲<'�7)��M:/���6}�T(5We:QL	J�?�B��u�\�r�.&f�ǭM�G�sI�N�l�/KS�������jn)Y8If�����q/D ?���H�N�G�e��r��6K�%Șvv�M|���vH�B~���"j��l���l�5����#�(�i���yP��Z������s�1n6�M�>P^<-��K�vѧ�c+�){�q�Y��8�=V;�!g���
�V��6-�aA��(�׵�J��(�K�Th�)��"x�/{����8K�Y��`Ax��Y�O�I�0"2�K6m۽��B����u!��O�����%d�@T}TV�}[�dL3#H���6#4O��zxp�`Qh�}C���q��J����%���+*���I
����&�t%@�*6��ٝ.��l�	����e7� �:�~����'b�q:���S��1�l��s���ZcL4�p�'>����e9�[U"�xj1裵����
Od>G�f�\��J�s�S�ۇ[�·�����=�a��X�*rIp@��2�p�N��X�b1C��	�Ps ����׫C]�-�믠��B���g�۷�)��&j_(ìX�]/ٷ}`7P�L������ȩ����K�X	,�\#vO��\0Lw'�58ʔ��X�!���ϝ�����:8�����mJ�d �2k(�|Ku�d$-��݈a)���4�x������}��D��3q����E�����k�D[�K����q�����eV�κJ$3��Ew�������ҮA�ƅDf�;�_�@��T��+�F��Ibv*J��[�k��[���L��X�p��6kK6#�~dV�N^l���˧��f���د�����;�6�`�]�/�*�ps���9�����ۼQ BV������Ob~\���HxV_����,N�Vx{
F��5N*xQ|[�X�t����e`҅%��GƼµK�J��T��^b�r�Iȱu~��O�Q�I��C�7�q9�����T�������BV���zD�ju���;^j�BRT��_�*<��T�j��(�8�S��Q����bvN��}�Ozw�������D)�F�13��<��z�{8���R�u)�� <-�CA%��'�RY��Qg��l�I>4����S'��;�yҍ&�)�T����[N:�boǂ7���+�B��5���E�P	�\hJ��j�W�羁�A0��'u/Ϧ)�v��	�o���Рq%E�l��6D���G�� � � #oF���P�ؗ����$���kCDM��3�8!�f+�e��I@Z�3���a�h���w!�@YZ\{�Vk��t66+�6E�����v������%u?���X������c��p�^���� ���՗�Q�3S1����@�IÖ�������;p����`9�����i8�JѲ��zJ,����W̞*I� %d�[�l�-�e��(��o1z���?�bE��ކ/:�3)�1H�ag_��!	(��J�$���9ѩB������ ��5��.Gi���m�����Կ	ͅ��v9�£��,�N"	�'>�d�hb�D�I/:��x�o�q��J=D�2Ҁ�����*��X������̹|7��ס���]Ybk��q*j-2���owUD��q@�VP�fdF;_�˳Vjzq��Xم��}
yI�D��萻sqJ�6޺��2�(�⍴P����)	z�6�M$��Bu4%	f}}֢��rQ��}�;[9%Ӹ(��������/��A��$�bx8G*^�2��h�6����P��2�/��M�R�V^��M�S���M�f@��Jz�̑ ���,���-�;1�?
͒�QC�(k�{'i�����؟�
�=��;��
�C���HN���f��Rz�3��?����b�U�Թ�Z�5��H�ܩ�[+���u��q�qT��`�QYv6��܏gu��lQ9U��l}+o�%;]�WbH���}��M�!�#�����l^�	�}�q޿�5�@��{v���կA�T�5����O�&c��O���]gd��F�xLҏ��2��(�Қ;��f�F-e祆�0:1�.�������;f�+�B�.����>#Q�����e!.Y��6���
��>:�%��$|W�l� P)�ȧ�c�8H�?sؠ#���VX7��}�3�8|�`��H0���%ʮn�~�E���*���"ȉ�������F�UʲYu�ـ�{�`\`�g����XHK��2�e�8ek0��y7H��'3�U���z�rY���GF&E������r+��k��a����^לp⨝��A�&��g��9�[X���8�!z��H�Y�:��P
8�#l=��M��1�*�/�u�r����6#oxBDI��xs��[ș�׊:�RE.J�� ��"��jv�d�Y��s�����6x8��g�t�"�#r-�����`,bB��T����]��,C���9��u=L@�a9�e�S�?���Ln�O���� $v�=Ӭ�p^$<�*?�C�j����q`�1{=�9�ϸ�����B��̣a5�4��>QޞX��:2`�$���I��M_KNn~n*a]�2/g8@�	C��δ�^��MM���B����H,e]����	��a1[��auK��t���G:��c�(e+���Ӈ*P�怼j��bTަ_l/�b��U�)�D�=�܏�ە;����<��ߠ��H�ә)�{
�βi)�+*we�g�:u�?l��Iǝ�A�@��Y�*�W'�y,��~R�m&[}+�1�4y����$gg���r�9�&k�3V�c��3�}+hIs��CT+�ìv�-�'{
[|�Ӻʄ\I��K���t0
�(=��~����d]`)��%P��d�Q��� ,���l�6`b�67����I����W97������Q����k���h_����E��WY�C�|�?����ʁ�}��M�`�Q�����	n��רN�~hKG,��� �R^=,�\%��d5בT!�e��fD��U
����lE�_oU��������̍�s�%rAt��;�a�wɦ����x�o9���󃳼nNnP�cs����B�ޑ
;W�a]3�?n��8t�蓾�V��֮�}�u���<�e�]TS)C�,P��NyJh�AO/*��ϱ֔�o�I���}���\�+íQ8�-�B��tI�i.�xOOq��}��+ 맜jkk��¨J���?��Cz�������W�u�Nz����<9�4��Zb�R��i�q�!w���
� ��/)J5�f#�6�}^?����U�p���}p���VQ�T8���j�&~m��_&�r��4W����LK��?�!G*=����2�|EB*���Pђ��!aaM���HưsO�'������`Y!2����&]�6
��5V9��b)Ses��^�	1�2_�LIև�i�ˬ:0\y	���hG+��2+>D���L�{���`{{e�I�-��c�K�J�h�����h���K㨇�%r��ڬ�X��ve��R�,!��Q���g�qLg�N0ظ
�&���I6�h�k��c�`���{��#z�&���þPo���: ��^�X�6W�6U7��j
��5֛M>���)a��-���g��9�dd:����y���dD���\՚�@�6k4�0w��3��d������)�F�k����J
+���2�ܢ[��ׄm���#z���+E�}WĴ���Y�Q`~����f��LD������ii�j��goH|[�������d���&�`eL�n9�7�<l>`G�;x��~�>�쓉p�������t|���!�웎M��*�x���0OM��_]�+�$������ջ�aS�Y9�?�P`�j��ޓM����Y�q7�8����ƹ*��2�!ѳ
�UV&�7�A���#H����s�EB��4�5����O�`�H��F[D'|$�F��Ooя���%����!g-Q�tɬ�1���o��L���O��q_���p��h>���h�-�,bZ)�=�~��0�P��s��P�C�ڋ��o����Ġ�� ��A΅"���5�3+����D1��!��i�m>��e�,�����]M.�W�� ��%�Pm6��yu]���g$d�|$�k +�R�;�-��$�S0�ZJ��Z��#�̸���F��y{��� �jE�N���=99p��Ъ�K;/�4LnC�B����v�������,2�O6�ˌ�HC�>?kQ�=��Lu�	:Ǫauv��0�ۚ݇|F�-ǔ�Zj�8^�&O�/n�k��N���f��%Y�#�Y�E���N�^&`�Я"���[�*�"�-�����3}GG�t��͵��2{6��ҙ��a�l�� .[�,��`��ɢV�x�;�GG�1I���[(��o�C�I�ڢ�%��Ȅ��l���+)���P�]Sz�$8�A�G>[.j�[�T��ꏼP#���y´�iN�b�&�[ʈ�q���6&�c�J��(a4��f�F?�Ճ��B�y��e�C��\-��%�s]�i��_�5 mMI�GЄ�8|�������"��S��4 ��M�����uć'M�)pn��{�s�X�*]�@�D���A�.�2���1��}�,i~g������qǇb�Q׶�7Iiu_��4$;���M�<�n6�0f��x�~-z���wD����p�G/o���R��=�ATXӡvg�B�fq�?�g��*t��**C�\Bd|��9����_�w�%�3��N~6��Y4,�9#�����/A�2͘��.����^��� [����,��i�yG��aR�x�]�S��G�5��I�Ӟ���!��U#�ƚ�ETI~P錨���2D�N�:ZM�6�R�	����M��i
��	7XwKZЏ�����WRCL_�V����[5�
�%j��������r+!�.����
`[p�qo&��}��M�x+X�2�+�*�hBf�YW�;�<���0gO&o�J�rURi�9�Aܾ{#o�Qf��T �	Ip^>//,�rM�,��Q�'O��7U����+�SJ���5�;߆��N��] ���;�C�a�Dj��u��*�(�+Q����Q_�Qmh�$Tt�s�X��s[�1m#[�s�,o���=YVg�����|.Q0ܯ���!��ߒ����v��H�MZ'"�|�c0��z�Z;�\��{��2S試܄�WOm�Q�:�x��ӆ�P]�@���֩MUd��ϻM��G��������,�*J�����%�I��M�'�Hڇ�*ӌn`l-2>߶�j�i���TZ��)z��d{t�R����N�{N|r����ۼ��^mt�hx�`%���10�Q[u7a��n�B�M��:1�E'98=�ϏM� ���[L#z���m� d�ڔ�-$aF�P��b�9�Y)�v���|Ǣ��Ch�2{7�p�(Q*^6��#��$�˘�����$��C�d�VP"��
=mQ�ie��4��Y�=Wa������͇�#��Y���c�_�<f��͋+}�A��%H����gO��������G����Z[����?��;~�i���6B��,]�f4t=\�z�^@ӀPށ�R,Q¡�ϼa
�Xy6�9ȀɰJv�2:��bf�6 ���x<Ki|im��#
.3�����yz��,]#0��p�<��\f ��7I6��.�B ��&�3�D��$D�������%,:	kq���r;�Hw�H4��r)in��I���&B�>�F^w"n��h���R��ͨv	�YRX#�.|���藧��X�S/L�H�1ږ�W�R]+Wa� �=
O���YG7��Ξ=J�h"*GLV��?��sǹ