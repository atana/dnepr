XlxV38EB     8f8     1ff:�&�S�Pn8beٍJz��L'�xN<��J���z���sp�z��Ի�뫑����jp�m2���(��C�e9k�!�P��ek�	r��2��q}?$�
��xW�������j�O3~SrK~���
v�Nbx�,H̱%^��i��w�_����O%)�Ւ�l@Ջ�%��d�����E&ȿ��� 	e�捊ݟ��I�B������r�����L���ަ���0����I�G��Ei�M�G�PZ�]_�G�̀"�	������hI)LS��j��
W*@T}D�Swd����������2Û�nD���#����Y�B0ub�β�}��f.���<�ٲ��,�d�=}��� z�L�X\:���r ۧ��`0k-&���`>PF"�-��)"GBh�샏ىe�6�y������ ����N-�Lǃ^9��ʅF��֮>�}��H�A+D�K��>Q��k~�	���S�ٞz�>���ۓ�)ȫ�,�6o֩�!f�j�N��2fs