XlxV38EB    1678     5caȜwJ=]Ã�h��gtP����ܩ�lj�L�2�������z���  N�IX�&��ʪ݊��� +�e����"4P����,<���5V=�Q�;q�	��[�
Oh��?sM��"^����ҔAz�b<z�g���m�QAL=v[�!_��'< 䖰�# I*ߎ
��ؓ>�4`�#�x��"m�	c䙕x��\W[(�K_�v����<��/t2G�H��#�Ԑ�P��ڍ��)`e��j1$u{�n�q������('�*�@���6+��r[�j�`�>��D�h&m0h�2��|�-��3j�C�jZO��X��ߵ�_��TD-�j�y_�ֳ��;
��<��kUVs�x�"��n
�.�E���a��B$���n\-�22��{�R�i;Rd������D&O���V������P��2:��G�7s��'xc��Z����O(l����g�p����`ys�"WE�c����ܵ��wQ������[>�c^~�%�<VXs������:!Q��,;��\�fu�	X�N�7�M��������x��g�/����X����0Q\���� �͂EM���ӥ�~[���y7xV�H#}˙H�ML�yE� ������똴��$<�L�Z�Ǧ(���.�+���?�m~�%F����� dnXO�bA��0\E$��"+)��K/)@k����O��n�7z��!����`���&�]v=D�G��$8K;�}ҟ�g{d`^gU8�ΔG&˛��-��������J���s{<�W���0�s�$*���G9@����.��f%�E�|8G2�.Vj����O��������.���C�5�5x�4��R�^ĀB�B'Zxk�[��f���ӿa�}�,������Y���K}nG?��=3	� �C���D�y���^�w�H����dPW�V�nA������	�-�d�����
�=fU�<.��>�Û��CG��f�%�C̢%O�>�F�#�c9tZ��7�/$оmܹ:I�����M�9����ӏ��5�-(<�2���G��%^ǝ�#�" ��6��K����qC}�u��m/<7��,�|8�*����#cO�G�76'8���=�G�Rm��uj�t��`�֢x��|'
�k���]�Z�V��3��"�=mv0H�V��\��hV��-^�QI�i;楥�k�����%��d��[��c��ڭ���m�4[B��f�L�E�E���:ПO�*��f��h�u{@y�B�cF���:Vȧ@|���Yy�劓�e>��L^߾0�*���~�q�c^����k���H�N��e����#Ŭ���4��"L��3���D~���4_�4F�N��jvN�E>�����H*Ø��y�Q�6�pu����=Bb�A(�\��S�L��xܥ�EY���I�)c)8,!�xߴ@Li�v�l�{�