XlxV38EB    12e1     4c6��A�� >�D��I"���z·���~Ӿ�9*�Z2�^G��$q/����{�h@>�+��i�-j4G��v�y���a�.��DtX�:���g����mp&��̩Y�`T���h�T.��:��E�\��cZ@J���)�_�1_�UU�J}(1�8q �S�&���!��tF-���=�sH������dp }'��~�m��	[W~{�����<K�
0+_����2vI�d���0a!�?�����Ә��� �xP�R��-4u�JC�5������Z�_-s�L��a@S��1t{��n}�����z'�$M��@�u.�}�x�1N�o	wrZɩR��A�{��`O��Uq�ݽ�$=����D
0��'D�z��f�����(�ڭ���i}¤=��t�n�˒9Dl���|�V;��Y�t���gϱשD����΃�&laX�̋g�P�Y0�PߞI�A���6��{����n��2�2O�v����d����#}��b��7.*��,q����}�(��;:��t�J(��4�� U�bӥ����m@y�#]]�M��:���<p��� C\*�I�Ħ���~����˯�Ken1���4��r��#��d�"1h���bD7fH"6> �#�6��u�=�IѢ� �]IԘ[o�U�d��j]&`��b5d�|��I��A��!��"jޗ������*�8|��\<{U5md\��3�țP�;2�dj2>�<�%�V8D���]e��j4F�x��4C���Z�t"�6x�'D� �"!�?�G~��q�8O����.�u���>�q��kB6oē�`�c8{���7Ă;T\�W�)R"�#������2�����=X�������F3�:�"(�����.��R[r�+����6�T�Z�EQ��؟j^!uE��Չ}wO.�(/��,�V�SWgÜ�~�LzD.Jc�
��ݲ����"���)���� 1��{�W��@�҆���ȧ���PpNYv�\���V\���x3(�h��r��"}��'�5ܚs�t����L��}���ďF��W��cv����Q�����1;�
��1�������� U��������n|G�ljg+��Qʅ=#�v{�Q|-D���l�R�B��bV�qKL0���r	<b�6pg���+��o�G\�.D�:rJ�@�@^�d�R�fk�~{���ń��1}H�a<�z�r