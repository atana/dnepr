XlxV38EB    1505     510}��_i�7�3��3m��۸fPͤ�B4� ���$[�����{:�g灶��c����1?����.��Ҵ��� ��B�C����{�U-ʡ̉���'��$5��+�'4l(:�j�I����r��NTm#�xY�ĉ�S��,����K��w1��5GȬMT���)�c�ֻ�hv��s,���q�f4-�䅞���K/�:ɈQ��,
��X��4��%x^��;J��f��+�ԋR��fk�l�U���/�@�!&�as���&�B��e'x ��4w�g�R����'6��H� ����hxv�� �DB�	^*eC7�j�t��̲Yn%CdV�֮i��&���|W�h�师��:����m�2���N��CBǼ��6�n_zš2b\\�&�\�=ѫ�ʛ�g�:^I����|1)o�X`m�9k�e�o�������ǮK�E5��'noL
�'�569�R���Y�ᥝ��dH�h������V<hd���w����Ә���2�A�~� �j��Zh[/��2�)����;�N����揋�Z��i�+a��`�Z��8'X	s���������g������6�T�Kji����������z�t��e�t�V���L��r��&���^��.��5�R�lp�M}<L�!��d��W��;;46�:=������bl`�|ss%�!���d`��G��qC��y�e�d^�)k�[�h� Ŝ�b���5���R�`�O �+�++��3�v9�O3-��d�>В>b�]�؞?�n�5��ڣ�-@,�))St[-.�����T)��Wů�Ȇ�.�~@g��� ���G���|�ߍ���w��>�g��g*j̓vQ���M�� c��4�T-��CAb�z�� z�Ȳ�ŢH�~qf��4{��D5H Mݿw�;	�Y�e;̯r>�ɡ�� ��?٭.0H�?�c�ad`E��RW�P�����OC�M&a����Z�^�V7��,�=�u>�_� ��<d2�=aL�1�.��=d&8"�]S1��f+;!z& �P0��r�b���r�r�k�lt糡�c�0��Z��G�W���>�g��t�7�p�
ܸ�x��C K���B�BP��:���\p�$�iG�P�=<!V�!#�����޺�%fڋR��߳�Y��j\ߞv~>*=p�Tvk�h�c��"T�n���C�N�)I���A�y�`��L���9�BE�5fpl�]�$�����ޠ���Q۲$7��_ a ���R��2