XlxV38EB    1366     4fc�6j�-{`%�J�<3s]f�7�,���ʌ��t�	���$ҧim�|�--c�8H��%�ޱ|f�LG���I��xbK*W�Zu��y�;t]vd�?��ك�Ȳ��M~V���|�J�upȦ,��R���|�!x�.Ī�k��9���V�tĊ��ĵ���#�t�b:��|)���^�G�
�;>w?$A���a�'��.q�d
O�W��R1�0H?���Q�SC��q ��ӻ�>����H[�t��:Q#��؋r�F�ҍ)��^�G+��Kr>{+�KLZ>�A���3(m�_>E�N��4�\5Q�˷�����@��oTM͹!}*���7�.!!�l��n�$���(��I4~�GPZ�O����Ӽ�0<�N�eo�����K�7����K�C�{���(�UJ�"$���a�犄B�hx�y�q��w mJ��B����`�i�h)^@ע�lfpa�n����2�|������s)�7疮�Vy�����&�rQ}�K )8�]��i��`�����J� rr�vhI��;b�R�e�����eN���^I�]7pΗ7��r曹��v�6�%��c����G��ј2f��qd[��� .[$ߺ5�K0�8Gc���L����d��b.\�?�Ş��l,C�6縼��b�ѝmB�rCj��������21�}�l�Nro�I���h>��͂�p�Ĺ����G���'���ѧ�y�$�Z3�R;D�9!_XW�'������X�Vw+)��r���Z��{OOL@"���Σ�x�	���ʮ�����ً7B̙:�ӧ��t�.FB\3�}/�����m/����l'���Љ:
����㫞�8�L��T2,���2�7�<s�?)��q�uh'X���T���L/_�o�p�:r�~*�(o�Q$�6sp��$�U�g<w���=�{�Cb�s��{�|�f=���G �QE�bU�c@����5���ޣ^j��u���d�\��yKanml3LN��C�6ò�.I����t��{-H��P8V��O���l��4�PNM�簉��]G�<!vz�y@7���L��or�j߰�ym>D�K�e*D�o՝>`�i���IN�-И[��Fa�-$��)��E���d���ģvePʵ�����X��#�F��lB&׋�D0��zCvA��k(��`�Ym"�r�P �^ʊ�ҧBUcOH,>؏�Pۖ��+���[�#�,�)m�;PA�O_r3pf��)�ftV���'K�U�P